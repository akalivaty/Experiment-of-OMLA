//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n212), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n222), .A2(G97), .ZN(new_n245));
  INV_X1    g0045(.A(G97), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n229), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n203), .A2(G20), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n253), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n207), .A2(G1), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G50), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G50), .B2(new_n263), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT66), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(G226), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G222), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G223), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n274), .C1(G77), .C2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n289), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(KEYINPUT9), .B2(new_n270), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n270), .B1(new_n296), .B2(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n282), .A2(new_n298), .A3(new_n288), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n277), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n281), .A2(G238), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(G232), .A4(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT67), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n283), .A2(KEYINPUT67), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(G226), .A3(new_n285), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n274), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT13), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n306), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n322), .C2(new_n296), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n305), .B1(new_n274), .B2(new_n316), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT68), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n318), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n329), .B2(new_n318), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n331), .A3(G179), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n296), .B1(new_n319), .B2(new_n321), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n323), .A2(new_n332), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n259), .A2(G77), .ZN(new_n339));
  INV_X1    g0139(.A(G50), .ZN(new_n340));
  INV_X1    g0140(.A(new_n260), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n339), .B1(new_n207), .B2(G68), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n264), .A2(new_n214), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n265), .A2(G68), .A3(new_n267), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT11), .B1(new_n342), .B2(new_n253), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT13), .B1(new_n326), .B2(KEYINPUT68), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n318), .A2(new_n329), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n325), .B(new_n327), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n352), .B1(new_n355), .B2(new_n291), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT70), .A4(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n349), .B1(new_n322), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n254), .A2(new_n263), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n256), .A2(new_n266), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(KEYINPUT75), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n365), .A2(KEYINPUT75), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n264), .B2(new_n256), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT73), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n308), .A3(G33), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n308), .B2(G33), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n258), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n207), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n207), .C1(new_n373), .C2(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(G68), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n214), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n202), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n260), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n254), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n283), .B2(G20), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n307), .A2(new_n309), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n207), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n214), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n388), .B1(new_n396), .B2(new_n387), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n369), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n370), .A2(new_n372), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  INV_X1    g0200(.A(G226), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n399), .A2(new_n402), .A3(new_n375), .A4(new_n376), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n274), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n277), .B1(G232), .B2(new_n281), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(G179), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n274), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n403), .B2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n281), .A2(G232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n303), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT18), .B1(new_n398), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n381), .A2(G68), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n375), .A2(new_n376), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n399), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n380), .B1(new_n419), .B2(new_n207), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n389), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n253), .A3(new_n397), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n368), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n414), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n406), .A2(new_n291), .A3(new_n407), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n359), .B1(new_n410), .B2(new_n412), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n428), .A3(new_n368), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n422), .A2(new_n428), .A3(KEYINPUT17), .A4(new_n368), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n416), .A2(new_n425), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n265), .A2(G77), .A3(new_n267), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n256), .A2(new_n341), .B1(new_n207), .B2(new_n220), .ZN(new_n435));
  XOR2_X1   g0235(.A(KEYINPUT15), .B(G87), .Z(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n259), .B2(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n434), .B1(G77), .B2(new_n263), .C1(new_n437), .C2(new_n254), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n283), .A2(G238), .A3(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n283), .A2(G232), .A3(new_n285), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n222), .C2(new_n283), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n274), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n277), .B1(G244), .B2(new_n281), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n438), .B1(G190), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n359), .B2(new_n445), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n296), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n438), .C1(G179), .C2(new_n444), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR4_X1   g0250(.A1(new_n302), .A2(new_n363), .A3(new_n433), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n264), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n254), .B(new_n263), .C1(G1), .C2(new_n258), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n454), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n207), .C1(G33), .C2(new_n246), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(G20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n253), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT20), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n457), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT21), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n469), .A3(new_n296), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n418), .A2(G264), .A3(G1698), .A4(new_n399), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n393), .A2(G303), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n418), .A2(G257), .A3(new_n285), .A4(new_n399), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n373), .A2(new_n377), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT78), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(G257), .A4(new_n285), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT79), .A3(new_n474), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n409), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n279), .A2(G1), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n274), .A2(new_n275), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G270), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n409), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n470), .B1(new_n487), .B2(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n479), .B(new_n473), .C1(new_n483), .C2(new_n484), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT79), .B1(new_n485), .B2(new_n474), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n274), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n468), .A2(new_n298), .A3(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n466), .A2(new_n467), .ZN(new_n503));
  INV_X1    g0303(.A(new_n457), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G169), .ZN(new_n506));
  INV_X1    g0306(.A(new_n496), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n497), .B(new_n502), .C1(new_n508), .C2(KEYINPUT21), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n500), .A2(G190), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n480), .A2(new_n486), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n496), .B1(new_n512), .B2(new_n274), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n511), .B(new_n468), .C1(new_n513), .C2(new_n359), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n453), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n469), .B1(new_n513), .B2(new_n506), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n500), .A2(new_n507), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n470), .B1(new_n500), .B2(new_n501), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n518), .A4(new_n453), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G250), .A2(G1698), .ZN(new_n522));
  INV_X1    g0322(.A(G257), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n418), .A2(new_n399), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n495), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n274), .B1(new_n528), .B2(G264), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n493), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n298), .B2(new_n530), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT23), .B1(new_n222), .B2(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n534), .A2(new_n535), .B1(G20), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n283), .A2(new_n207), .A3(G87), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n538), .A2(new_n216), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n418), .A2(new_n207), .A3(new_n399), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n540), .B2(new_n543), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(new_n254), .ZN(new_n546));
  OR3_X1    g0346(.A1(new_n263), .A2(KEYINPUT25), .A3(G107), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT25), .B1(new_n263), .B2(G107), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n456), .C2(new_n222), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT83), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n533), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n545), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n253), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n549), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT84), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n532), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n530), .A2(G200), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n529), .A2(G190), .A3(new_n493), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(new_n554), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n493), .B1(new_n523), .B2(new_n495), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n399), .A2(new_n285), .A3(new_n375), .A4(new_n376), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n221), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(new_n458), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n563), .B1(new_n570), .B2(new_n274), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n298), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n246), .A2(new_n222), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n573), .B2(new_n245), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n392), .A2(new_n395), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G107), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n253), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n264), .A2(new_n246), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n456), .B2(new_n246), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n572), .B(new_n586), .C1(G169), .C2(new_n571), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n571), .A2(G190), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n584), .B1(new_n581), .B2(new_n253), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n571), .C2(new_n359), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n215), .A2(new_n285), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n221), .A2(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n418), .A2(new_n399), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n409), .B1(new_n594), .B2(new_n536), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n409), .B(G250), .C1(G1), .C2(new_n279), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n492), .A2(new_n489), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n456), .A2(new_n216), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n601), .B(KEYINPUT77), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT19), .B1(new_n259), .B2(G97), .ZN(new_n603));
  OR2_X1    g0403(.A1(KEYINPUT76), .A2(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT76), .A2(G87), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n575), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT19), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n314), .B2(new_n207), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n418), .A2(new_n207), .A3(new_n399), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n214), .ZN(new_n611));
  INV_X1    g0411(.A(new_n436), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n253), .B1(new_n264), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(G200), .B1(new_n595), .B2(new_n598), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n600), .A2(new_n602), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n456), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n599), .A2(new_n298), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n296), .B1(new_n595), .B2(new_n598), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n591), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n452), .A2(new_n521), .A3(new_n562), .A4(new_n623), .ZN(G372));
  AOI21_X1  g0424(.A(new_n360), .B1(new_n356), .B2(new_n357), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n351), .B1(new_n625), .B2(new_n449), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n431), .A2(new_n432), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  AOI221_X4 g0429(.A(KEYINPUT18), .B1(new_n413), .B2(new_n408), .C1(new_n422), .C2(new_n368), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n424), .B1(new_n423), .B2(new_n414), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n416), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n300), .B1(new_n635), .B2(new_n295), .ZN(new_n636));
  INV_X1    g0436(.A(new_n561), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n591), .A2(new_n637), .A3(new_n621), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n554), .A2(new_n556), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n532), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n509), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n638), .B(KEYINPUT85), .C1(new_n509), .C2(new_n640), .ZN(new_n644));
  INV_X1    g0444(.A(new_n587), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n615), .A2(new_n620), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT26), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n621), .A2(new_n587), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n620), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n643), .A2(new_n644), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n636), .B1(new_n452), .B2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n551), .A2(new_n557), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n558), .A2(new_n661), .A3(new_n561), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n558), .A2(new_n661), .A3(KEYINPUT87), .A4(new_n561), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n558), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n660), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n660), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n468), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n487), .A2(new_n291), .A3(new_n496), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n359), .B1(new_n500), .B2(new_n507), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(new_n505), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT81), .B1(new_n674), .B2(new_n509), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n675), .B2(new_n519), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n509), .A2(new_n671), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n669), .B(G330), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n640), .A2(new_n670), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n664), .A2(new_n509), .A3(new_n670), .A4(new_n665), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n210), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n606), .A2(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n228), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n622), .A2(new_n558), .A3(new_n561), .A4(new_n670), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n515), .B2(new_n520), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n529), .A2(new_n493), .ZN(new_n694));
  NOR4_X1   g0494(.A1(new_n694), .A2(new_n571), .A3(G179), .A4(new_n599), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n517), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n496), .A2(new_n298), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(new_n599), .A3(new_n529), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n571), .A4(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n571), .A2(new_n697), .A3(new_n529), .A4(new_n599), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n487), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n660), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n690), .B1(new_n693), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n652), .A2(new_n670), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n638), .B1(new_n509), .B2(new_n667), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n620), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n649), .B2(KEYINPUT88), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT26), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT88), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n648), .B1(new_n621), .B2(new_n587), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT29), .B(new_n670), .C1(new_n714), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n709), .B1(new_n712), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n689), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n206), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n683), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n676), .A2(new_n677), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(G330), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n730), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n229), .B1(G20), .B2(new_n296), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n207), .A2(new_n291), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n298), .A2(G200), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT90), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT90), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(G190), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT92), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(KEYINPUT92), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n740), .A2(G322), .B1(new_n746), .B2(G329), .ZN(new_n747));
  NAND3_X1  g0547(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n291), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n207), .B1(new_n743), .B2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n748), .A2(G190), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n741), .A2(new_n736), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n359), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n735), .A2(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n393), .B1(new_n758), .B2(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n742), .A2(new_n744), .A3(new_n761), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n763), .B1(G283), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n747), .A2(new_n757), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n758), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n740), .A2(G58), .B1(G77), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT91), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n745), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n762), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n604), .A2(new_n605), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n393), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n755), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n778), .B2(new_n214), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n750), .A2(new_n340), .B1(new_n752), .B2(new_n246), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n774), .B(new_n781), .C1(new_n222), .C2(new_n764), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n767), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT94), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n734), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  INV_X1    g0586(.A(new_n729), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n682), .A2(new_n393), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n788), .A2(G355), .B1(new_n454), .B2(new_n682), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n481), .A2(new_n682), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n687), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n244), .A2(new_n279), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n207), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n734), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT89), .Z(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n787), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n795), .B(KEYINPUT95), .Z(new_n800));
  OAI211_X1 g0600(.A(new_n786), .B(new_n799), .C1(new_n730), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n732), .A2(new_n801), .ZN(G396));
  INV_X1    g0602(.A(KEYINPUT100), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n447), .A2(new_n449), .A3(new_n670), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n650), .B1(new_n641), .B2(new_n642), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n644), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n438), .A2(new_n660), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n447), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n449), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n449), .A2(new_n660), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n806), .B1(new_n710), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n787), .B1(new_n812), .B2(new_n709), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT99), .ZN(new_n814));
  INV_X1    g0614(.A(new_n804), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n652), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n660), .B1(new_n805), .B2(new_n644), .ZN(new_n817));
  INV_X1    g0617(.A(new_n811), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n693), .A2(new_n708), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G330), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n814), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n812), .A2(KEYINPUT99), .A3(new_n709), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n733), .A2(new_n794), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n729), .B1(new_n826), .B2(G77), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT96), .Z(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n216), .A2(new_n764), .B1(new_n745), .B2(new_n759), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G294), .B2(new_n740), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n778), .A2(new_n832), .B1(new_n758), .B2(new_n454), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT97), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT97), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n752), .A2(new_n246), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n393), .B1(new_n762), .B2(new_n222), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G303), .C2(new_n749), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n481), .B1(new_n340), .B2(new_n762), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n214), .A2(new_n764), .B1(new_n745), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n752), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n840), .B(new_n842), .C1(G58), .C2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT98), .Z(new_n845));
  AOI22_X1  g0645(.A1(new_n768), .A2(G159), .B1(G137), .B2(new_n749), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n778), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G143), .B2(new_n740), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT34), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n839), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n829), .B1(new_n851), .B2(new_n733), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n818), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n803), .B1(new_n824), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n822), .A2(new_n823), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT100), .B(new_n854), .C1(new_n857), .C2(new_n813), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n726), .A2(new_n206), .ZN(new_n860));
  XOR2_X1   g0660(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n861));
  INV_X1    g0661(.A(new_n387), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n417), .B2(new_n420), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n388), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n369), .B1(new_n390), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n429), .B1(new_n865), .B2(new_n658), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n415), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n658), .B1(new_n422), .B2(new_n368), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n423), .A2(new_n414), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n429), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT16), .B1(new_n382), .B2(new_n862), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n421), .A2(new_n253), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n368), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n658), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n433), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n873), .B2(new_n880), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT103), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n876), .A2(new_n414), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n878), .A3(new_n429), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n871), .A2(new_n429), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(KEYINPUT37), .B1(new_n888), .B2(new_n870), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n630), .A2(new_n631), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n878), .B1(new_n890), .B2(new_n627), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n885), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n873), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n349), .A2(new_n670), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n351), .A2(new_n362), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n350), .B(new_n660), .C1(new_n625), .C2(new_n338), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n811), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n691), .B1(new_n675), .B2(new_n519), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n706), .A2(new_n707), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n861), .B1(new_n895), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n423), .A2(new_n877), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n871), .A2(new_n905), .A3(new_n429), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT104), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n869), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n634), .A2(new_n627), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n869), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n893), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n820), .A2(new_n912), .A3(KEYINPUT40), .A4(new_n900), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n451), .A3(new_n820), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(G330), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n451), .B2(new_n820), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT106), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n338), .A2(new_n350), .A3(new_n670), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n892), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n908), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n906), .A2(new_n908), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n431), .A2(new_n432), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n632), .B2(new_n633), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n924), .B(new_n925), .C1(new_n927), .C2(new_n905), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n881), .B1(new_n928), .B2(new_n885), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n922), .B(new_n923), .C1(new_n929), .C2(KEYINPUT39), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n632), .A2(new_n633), .A3(new_n658), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n898), .A2(new_n899), .ZN(new_n933));
  INV_X1    g0733(.A(new_n810), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n933), .B1(new_n806), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT102), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n895), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n933), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n816), .B2(new_n810), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT102), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n932), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n451), .B(new_n722), .C1(new_n817), .C2(KEYINPUT29), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n636), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n941), .B(new_n943), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n860), .B1(new_n920), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n920), .B2(new_n944), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(G116), .A3(new_n230), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n201), .A2(G68), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT101), .Z(new_n952));
  NOR3_X1   g0752(.A1(new_n687), .A2(new_n220), .A3(new_n384), .ZN(new_n953));
  OAI211_X1 g0753(.A(G1), .B(new_n725), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n950), .A3(new_n954), .ZN(G367));
  NAND2_X1  g0755(.A1(new_n645), .A2(new_n660), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n587), .B(new_n590), .C1(new_n589), .C2(new_n670), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n680), .A2(new_n679), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n679), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n680), .A2(new_n679), .ZN(new_n964));
  INV_X1    g0764(.A(new_n958), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT44), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n964), .A2(KEYINPUT44), .A3(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n678), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n666), .B(new_n668), .C1(new_n510), .C2(new_n660), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n680), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n730), .A2(G330), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n676), .A2(new_n677), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n680), .B(new_n971), .C1(new_n974), .C2(new_n690), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n963), .B(new_n678), .C1(new_n966), .C2(new_n967), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n970), .A2(new_n723), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n723), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n683), .B(KEYINPUT41), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT108), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT108), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n983), .B(new_n980), .C1(new_n978), .C2(new_n723), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n727), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n680), .A2(new_n965), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n587), .B1(new_n957), .B2(new_n558), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n670), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n670), .B1(new_n602), .B2(new_n613), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n715), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n621), .B2(new_n991), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n990), .A2(KEYINPUT43), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n993), .B(KEYINPUT43), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n990), .A2(KEYINPUT107), .A3(new_n995), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n994), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n678), .A2(new_n965), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n985), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n790), .A2(new_n240), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n798), .B(new_n1004), .C1(new_n210), .C2(new_n612), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT109), .Z(new_n1006));
  AOI22_X1  g0806(.A1(new_n740), .A2(G303), .B1(G311), .B2(new_n749), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT110), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n762), .A2(new_n1009), .A3(new_n454), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n762), .B2(new_n454), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n222), .B2(new_n752), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G294), .C2(new_n755), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n419), .B1(new_n832), .B2(new_n758), .C1(new_n745), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G97), .B2(new_n765), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1008), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n752), .A2(new_n214), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n283), .B1(new_n201), .B2(new_n758), .C1(new_n778), .C2(new_n771), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G143), .C2(new_n749), .ZN(new_n1020));
  INV_X1    g0820(.A(G137), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n745), .A2(new_n1021), .B1(new_n383), .B2(new_n762), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT111), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n764), .A2(new_n220), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n740), .B2(G150), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1017), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n787), .B(new_n1006), .C1(new_n1031), .C2(new_n733), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n800), .B2(new_n993), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT113), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1003), .A2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n976), .A2(new_n728), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n237), .A2(new_n279), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(new_n790), .B1(new_n686), .B2(new_n788), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n257), .A2(new_n340), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n279), .B1(new_n214), .B2(new_n220), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1041), .A2(new_n686), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1039), .A2(new_n1043), .B1(G107), .B2(new_n210), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n787), .B1(new_n1044), .B2(new_n798), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n740), .A2(G50), .B1(new_n746), .B2(G150), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n762), .A2(new_n220), .B1(new_n758), .B2(new_n214), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n419), .B(new_n1047), .C1(new_n765), .C2(G97), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n749), .A2(G159), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n612), .A2(new_n752), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n755), .B2(new_n257), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT114), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n768), .A2(G303), .B1(G311), .B2(new_n755), .ZN(new_n1054));
  INV_X1    g0854(.A(G322), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n740), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1054), .B1(new_n1055), .B2(new_n750), .C1(new_n1056), .C2(new_n1014), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n775), .A2(G294), .B1(new_n843), .B2(G283), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n419), .B1(new_n764), .B2(new_n454), .C1(new_n751), .C2(new_n745), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1063), .B2(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1053), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1045), .B1(new_n1067), .B2(new_n734), .C1(new_n669), .C2(new_n800), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n976), .A2(new_n723), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n683), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n976), .A2(new_n723), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1037), .B(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(G393));
  NAND3_X1  g0872(.A1(new_n970), .A2(new_n728), .A3(new_n977), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n790), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n798), .B1(new_n246), .B2(new_n210), .C1(new_n250), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n729), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n740), .A2(G311), .B1(G317), .B2(new_n749), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n393), .B1(new_n758), .B2(new_n753), .C1(new_n832), .C2(new_n762), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n778), .A2(new_n760), .B1(new_n752), .B2(new_n454), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n222), .B2(new_n764), .C1(new_n1055), .C2(new_n745), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n740), .A2(G159), .B1(G150), .B2(new_n749), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G87), .A2(new_n765), .B1(new_n746), .B2(G143), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n762), .A2(new_n214), .B1(new_n758), .B2(new_n256), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n419), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n752), .A2(new_n220), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n201), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n755), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1078), .A2(new_n1082), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1076), .B1(new_n1092), .B2(new_n733), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n958), .B2(new_n795), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n970), .A2(new_n977), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1069), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n978), .A2(new_n683), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1073), .B(new_n1094), .C1(new_n1097), .C2(new_n1098), .ZN(G390));
  OAI211_X1 g0899(.A(G330), .B(new_n818), .C1(new_n901), .C2(new_n902), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n938), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT39), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n912), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n935), .A2(new_n921), .B1(new_n1103), .B2(new_n923), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n912), .A2(new_n921), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n670), .B1(new_n714), .B2(new_n721), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n809), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n810), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n933), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n923), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n939), .B2(new_n922), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n721), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n660), .B1(new_n1113), .B2(new_n713), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n934), .B1(new_n1114), .B2(new_n809), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n912), .B(new_n921), .C1(new_n1115), .C2(new_n938), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n820), .A2(new_n933), .A3(G330), .A4(new_n818), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1110), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n709), .A2(new_n451), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n942), .A2(new_n1120), .A3(new_n636), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1100), .A2(new_n938), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1117), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1117), .A2(new_n1122), .B1(new_n816), .B2(new_n810), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n684), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1100), .A2(new_n938), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(new_n1101), .B1(new_n806), .B2(new_n934), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1117), .A2(new_n1122), .A3(new_n1115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n1110), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1110), .A2(new_n1118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n728), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1111), .A2(new_n794), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n729), .B1(new_n826), .B2(new_n257), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT115), .Z(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n283), .B1(new_n758), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n778), .A2(new_n1021), .B1(new_n750), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(G159), .C2(new_n843), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT53), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n762), .B2(new_n847), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n775), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n740), .A2(G132), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n746), .A2(G125), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n765), .A2(new_n1089), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1142), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n740), .A2(G116), .B1(new_n746), .B2(G294), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n750), .A2(new_n832), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1088), .B(new_n1151), .C1(G107), .C2(new_n755), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n393), .B1(new_n758), .B2(new_n246), .C1(new_n216), .C2(new_n762), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G68), .B2(new_n765), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT116), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n734), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1149), .A2(KEYINPUT116), .A3(new_n1155), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1137), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1135), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1132), .A2(new_n1134), .A3(new_n1160), .ZN(G378));
  NAND3_X1  g0961(.A1(new_n904), .A2(G330), .A3(new_n913), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n270), .A2(new_n658), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n302), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n302), .A2(new_n1165), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1166), .A3(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1162), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n904), .A2(new_n1172), .A3(G330), .A4(new_n913), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n941), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n941), .A3(new_n1175), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1131), .A2(new_n1121), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n683), .B(new_n1182), .C1(new_n1183), .C2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1173), .A2(new_n794), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n826), .A2(new_n1089), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n765), .A2(G58), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT117), .Z(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n778), .A2(new_n246), .B1(new_n750), .B2(new_n454), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1018), .B(new_n1190), .C1(new_n436), .C2(new_n768), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n740), .A2(G107), .B1(new_n746), .B2(G283), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT118), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n419), .A2(new_n278), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G77), .B2(new_n775), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1191), .B(new_n1192), .C1(new_n1193), .C2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1189), .B(new_n1196), .C1(new_n1193), .C2(new_n1195), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1194), .B(new_n340), .C1(G33), .C2(G41), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n762), .A2(new_n1138), .B1(new_n758), .B2(new_n1021), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G132), .B2(new_n755), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n843), .A2(G150), .B1(G125), .B2(new_n749), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n1056), .C2(new_n1140), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n765), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n787), .B(new_n1186), .C1(new_n1210), .C2(new_n733), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1180), .A2(new_n728), .B1(new_n1185), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1184), .A2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n1130), .A2(new_n728), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n729), .B1(new_n826), .B2(G68), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1050), .B1(new_n740), .B2(G283), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n393), .B1(new_n758), .B2(new_n222), .C1(new_n750), .C2(new_n753), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1219), .B(new_n1025), .C1(G116), .C2(new_n755), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n745), .A2(new_n760), .B1(new_n246), .B2(new_n762), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT120), .Z(new_n1223));
  OAI22_X1  g1023(.A1(new_n762), .A2(new_n771), .B1(new_n758), .B2(new_n847), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n419), .B(new_n1224), .C1(new_n746), .C2(G128), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n750), .A2(new_n841), .B1(new_n752), .B2(new_n340), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n778), .A2(new_n1138), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n740), .A2(G137), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1221), .A2(new_n1223), .B1(new_n1189), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1215), .B1(new_n1231), .B2(new_n733), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n933), .B2(new_n853), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1214), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n942), .A2(new_n1120), .A3(new_n636), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1128), .A2(new_n1236), .A3(new_n1129), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT119), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT119), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1128), .A2(new_n1239), .A3(new_n1236), .A4(new_n1129), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n981), .A3(new_n1125), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1235), .A2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(G375), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT122), .Z(new_n1245));
  AOI21_X1  g1045(.A(new_n1034), .B1(new_n985), .B2(new_n1002), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(G378), .A2(G390), .A3(G381), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(G407));
  OAI21_X1  g1048(.A(new_n1160), .B1(new_n1119), .B2(new_n727), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1131), .B2(new_n1126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n659), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G375), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT123), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1252), .B(new_n1253), .ZN(G409));
  XNOR2_X1  g1054(.A(G393), .B(G396), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1255), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n1259), .A3(G390), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G390), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1174), .A2(new_n941), .A3(new_n1175), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n941), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1236), .B1(new_n1133), .B2(new_n1130), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n683), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1212), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1180), .A2(new_n981), .A3(new_n1181), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n728), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1185), .A2(new_n1211), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1250), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1264), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n1236), .A4(new_n1129), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1280), .A2(new_n683), .ZN(new_n1281));
  AOI221_X4 g1081(.A(new_n1234), .B1(new_n856), .B2(new_n858), .C1(new_n1279), .C2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1235), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1277), .A2(KEYINPUT62), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT62), .B1(new_n1277), .B2(new_n1285), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1277), .A2(new_n1285), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1288), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1264), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1283), .A2(new_n1235), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1283), .A2(G384), .A3(new_n1235), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1264), .A2(G2897), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1300), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1292), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1262), .B1(new_n1289), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1290), .B2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1277), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1285), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1313), .B1(new_n1277), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1262), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1290), .A2(new_n1309), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1312), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1307), .A2(new_n1318), .ZN(G405));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1250), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1285), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1271), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G378), .B1(new_n1184), .B2(new_n1212), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1271), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1285), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1261), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1257), .A2(new_n1259), .A3(G390), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1320), .B1(new_n1327), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1262), .A2(KEYINPUT127), .A3(new_n1326), .A4(new_n1323), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(G402));
endmodule


