

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n766), .A2(n775), .ZN(n523) );
  AND2_X1 U556 ( .A1(n696), .A2(n686), .ZN(n685) );
  NAND2_X1 U557 ( .A1(n664), .A2(G8), .ZN(n671) );
  INV_X1 U558 ( .A(n664), .ZN(n647) );
  BUF_X1 U559 ( .A(n664), .Z(n674) );
  NAND2_X1 U560 ( .A1(n729), .A2(n731), .ZN(n664) );
  XNOR2_X1 U561 ( .A(n522), .B(n609), .ZN(n729) );
  NOR2_X1 U562 ( .A1(n553), .A2(n552), .ZN(n608) );
  NOR2_X1 U563 ( .A1(n590), .A2(n558), .ZN(n815) );
  BUF_X1 U564 ( .A(n541), .Z(n906) );
  INV_X1 U565 ( .A(n535), .ZN(n914) );
  XNOR2_X1 U566 ( .A(n543), .B(n542), .ZN(n545) );
  AND2_X1 U567 ( .A1(n533), .A2(G2104), .ZN(n541) );
  INV_X1 U568 ( .A(G2105), .ZN(n533) );
  NAND2_X1 U569 ( .A1(n608), .A2(G40), .ZN(n522) );
  INV_X1 U570 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U571 ( .A1(n746), .A2(n523), .ZN(n767) );
  NOR2_X1 U572 ( .A1(G651), .A2(n590), .ZN(n816) );
  NOR2_X1 U573 ( .A1(n682), .A2(n681), .ZN(n684) );
  INV_X1 U574 ( .A(G168), .ZN(n677) );
  XNOR2_X1 U575 ( .A(n676), .B(KEYINPUT30), .ZN(n678) );
  AND2_X1 U576 ( .A1(n694), .A2(n675), .ZN(n676) );
  AND2_X1 U577 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U578 ( .A(n534), .B(KEYINPUT17), .ZN(n547) );
  INV_X1 U579 ( .A(n547), .ZN(n535) );
  INV_X1 U580 ( .A(KEYINPUT23), .ZN(n542) );
  NOR2_X1 U581 ( .A1(n765), .A2(n772), .ZN(n766) );
  OR2_X1 U582 ( .A1(n698), .A2(n697), .ZN(n524) );
  NOR2_X1 U583 ( .A1(n671), .A2(n706), .ZN(n525) );
  AND2_X1 U584 ( .A1(n616), .A2(n615), .ZN(n526) );
  XNOR2_X1 U585 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n527) );
  BUF_X1 U586 ( .A(n608), .Z(G160) );
  INV_X1 U587 ( .A(n1001), .ZN(n703) );
  AND2_X1 U588 ( .A1(n678), .A2(n677), .ZN(n682) );
  INV_X1 U589 ( .A(KEYINPUT31), .ZN(n683) );
  INV_X1 U590 ( .A(G2104), .ZN(n532) );
  XNOR2_X1 U591 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n622) );
  XNOR2_X1 U592 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(G164) );
  AND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n908) );
  NAND2_X1 U595 ( .A1(G114), .A2(n908), .ZN(n530) );
  NOR2_X4 U596 ( .A1(G2104), .A2(n536), .ZN(n909) );
  NAND2_X1 U597 ( .A1(G126), .A2(n909), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT88), .B(n531), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U601 ( .A1(G138), .A2(n914), .ZN(n538) );
  NAND2_X1 U602 ( .A1(G102), .A2(n906), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(G101), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n909), .A2(G125), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT64), .ZN(n553) );
  INV_X1 U608 ( .A(KEYINPUT65), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n547), .A2(G137), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n908), .A2(G113), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X2 U613 ( .A1(G651), .A2(G543), .ZN(n811) );
  NAND2_X1 U614 ( .A1(n811), .A2(G89), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  XOR2_X1 U616 ( .A(G543), .B(KEYINPUT0), .Z(n590) );
  INV_X1 U617 ( .A(G651), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G76), .A2(n815), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT5), .ZN(n564) );
  NOR2_X1 U621 ( .A1(G543), .A2(n558), .ZN(n559) );
  XOR2_X2 U622 ( .A(KEYINPUT1), .B(n559), .Z(n812) );
  NAND2_X1 U623 ( .A1(G63), .A2(n812), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G51), .A2(n816), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U629 ( .A1(G64), .A2(n812), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G52), .A2(n816), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G90), .A2(n811), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G77), .A2(n815), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(G171) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G65), .A2(n812), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G53), .A2(n816), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT68), .B(n575), .Z(n579) );
  NAND2_X1 U642 ( .A1(G91), .A2(n811), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G78), .A2(n815), .ZN(n576) );
  AND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G299) );
  NAND2_X1 U646 ( .A1(G62), .A2(n812), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G50), .A2(n816), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(KEYINPUT81), .B(n582), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G88), .A2(n811), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G75), .A2(n815), .ZN(n583) );
  AND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G303) );
  INV_X1 U654 ( .A(G303), .ZN(G166) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G49), .A2(n816), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U659 ( .A1(n812), .A2(n589), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n590), .A2(G87), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G288) );
  NAND2_X1 U662 ( .A1(G48), .A2(n816), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT80), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G86), .A2(n811), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G61), .A2(n812), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n815), .A2(G73), .ZN(n596) );
  XOR2_X1 U668 ( .A(KEYINPUT2), .B(n596), .Z(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G305) );
  NAND2_X1 U671 ( .A1(G60), .A2(n812), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G47), .A2(n816), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G85), .A2(n811), .ZN(n603) );
  XOR2_X1 U675 ( .A(KEYINPUT66), .B(n603), .Z(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n815), .A2(G72), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(G290) );
  INV_X1 U679 ( .A(KEYINPUT90), .ZN(n609) );
  NOR2_X1 U680 ( .A1(G164), .A2(G1384), .ZN(n731) );
  NAND2_X1 U681 ( .A1(G1961), .A2(n674), .ZN(n612) );
  XOR2_X1 U682 ( .A(G2078), .B(KEYINPUT25), .Z(n979) );
  NAND2_X1 U683 ( .A1(n647), .A2(n979), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n679) );
  OR2_X1 U685 ( .A1(n679), .A2(G301), .ZN(n663) );
  INV_X1 U686 ( .A(G1341), .ZN(n993) );
  XOR2_X1 U687 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n629) );
  NAND2_X1 U688 ( .A1(n993), .A2(n629), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n613), .A2(n674), .ZN(n616) );
  XNOR2_X1 U690 ( .A(G1996), .B(KEYINPUT98), .ZN(n970) );
  AND2_X1 U691 ( .A1(n970), .A2(n647), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n614), .A2(n629), .ZN(n615) );
  XOR2_X1 U693 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n618) );
  NAND2_X1 U694 ( .A1(G56), .A2(n812), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n618), .B(n617), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n811), .A2(G81), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G68), .A2(n815), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT72), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G43), .A2(n816), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n994) );
  NOR2_X1 U704 ( .A1(n629), .A2(n970), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n994), .A2(n630), .ZN(n631) );
  AND2_X1 U706 ( .A1(n526), .A2(n631), .ZN(n645) );
  NAND2_X1 U707 ( .A1(n647), .A2(G2067), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G1348), .A2(n674), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n634), .B(KEYINPUT100), .ZN(n646) );
  NAND2_X1 U711 ( .A1(G66), .A2(n812), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT74), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G92), .A2(n811), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G54), .A2(n816), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G79), .A2(n815), .ZN(n638) );
  XNOR2_X1 U717 ( .A(KEYINPUT75), .B(n638), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X2 U720 ( .A(KEYINPUT15), .B(n643), .Z(n996) );
  NAND2_X1 U721 ( .A1(n646), .A2(n996), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n646), .A2(n996), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n647), .A2(G2072), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT27), .ZN(n650) );
  INV_X1 U726 ( .A(G1956), .ZN(n879) );
  NOR2_X1 U727 ( .A1(n879), .A2(n647), .ZN(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n655) );
  INV_X1 U729 ( .A(G299), .ZN(n825) );
  AND2_X1 U730 ( .A1(n655), .A2(n825), .ZN(n651) );
  NOR2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n653), .A2(n654), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n825), .A2(n655), .ZN(n657) );
  XNOR2_X1 U734 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U737 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n662), .A2(n663), .ZN(n696) );
  INV_X1 U740 ( .A(G8), .ZN(n670) );
  NOR2_X1 U741 ( .A1(G1971), .A2(n671), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT103), .B(n665), .ZN(n668) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n674), .ZN(n666) );
  NOR2_X1 U744 ( .A1(G166), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n669) );
  OR2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n686) );
  NOR2_X1 U747 ( .A1(G1966), .A2(n671), .ZN(n673) );
  INV_X1 U748 ( .A(KEYINPUT96), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n673), .B(n672), .ZN(n694) );
  NOR2_X1 U750 ( .A1(G2084), .A2(n674), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n670), .A2(n692), .ZN(n675) );
  NAND2_X1 U752 ( .A1(G301), .A2(n679), .ZN(n680) );
  XOR2_X1 U753 ( .A(KEYINPUT102), .B(n680), .Z(n681) );
  XNOR2_X1 U754 ( .A(n684), .B(n683), .ZN(n695) );
  NAND2_X1 U755 ( .A1(n685), .A2(n695), .ZN(n690) );
  INV_X1 U756 ( .A(n686), .ZN(n688) );
  AND2_X1 U757 ( .A1(G286), .A2(G8), .ZN(n687) );
  OR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(n527), .ZN(n699) );
  NAND2_X1 U761 ( .A1(G8), .A2(n692), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n698) );
  AND2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U764 ( .A1(n699), .A2(n524), .ZN(n716) );
  NOR2_X1 U765 ( .A1(G1971), .A2(G303), .ZN(n700) );
  XNOR2_X1 U766 ( .A(n700), .B(KEYINPUT105), .ZN(n702) );
  INV_X1 U767 ( .A(KEYINPUT33), .ZN(n701) );
  AND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  NAND2_X1 U770 ( .A1(n716), .A2(n705), .ZN(n708) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  INV_X1 U772 ( .A(n1002), .ZN(n706) );
  OR2_X1 U773 ( .A1(KEYINPUT33), .A2(n525), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U775 ( .A(n709), .B(KEYINPUT106), .ZN(n712) );
  NAND2_X1 U776 ( .A1(n1001), .A2(KEYINPUT33), .ZN(n710) );
  NOR2_X1 U777 ( .A1(n671), .A2(n710), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n714) );
  INV_X1 U779 ( .A(KEYINPUT107), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U781 ( .A(G1981), .B(G305), .Z(n1011) );
  NAND2_X1 U782 ( .A1(n715), .A2(n1011), .ZN(n722) );
  BUF_X1 U783 ( .A(n716), .Z(n719) );
  NOR2_X1 U784 ( .A1(G2090), .A2(G303), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G8), .A2(n717), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n720), .A2(n671), .ZN(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U789 ( .A(n723), .B(KEYINPUT108), .ZN(n727) );
  NOR2_X1 U790 ( .A1(G1981), .A2(G305), .ZN(n724) );
  XOR2_X1 U791 ( .A(n724), .B(KEYINPUT24), .Z(n725) );
  NOR2_X1 U792 ( .A1(n671), .A2(n725), .ZN(n726) );
  NOR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U794 ( .A(n728), .B(KEYINPUT109), .ZN(n746) );
  BUF_X1 U795 ( .A(n729), .Z(n730) );
  INV_X1 U796 ( .A(n730), .ZN(n732) );
  NOR2_X1 U797 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U798 ( .A(KEYINPUT91), .B(n733), .Z(n779) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n734) );
  XNOR2_X1 U800 ( .A(n734), .B(KEYINPUT92), .ZN(n777) );
  NAND2_X1 U801 ( .A1(G140), .A2(n914), .ZN(n736) );
  NAND2_X1 U802 ( .A1(G104), .A2(n906), .ZN(n735) );
  NAND2_X1 U803 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U804 ( .A(KEYINPUT34), .B(n737), .ZN(n744) );
  XNOR2_X1 U805 ( .A(KEYINPUT35), .B(KEYINPUT94), .ZN(n742) );
  NAND2_X1 U806 ( .A1(n909), .A2(G128), .ZN(n740) );
  NAND2_X1 U807 ( .A1(n908), .A2(G116), .ZN(n738) );
  XOR2_X1 U808 ( .A(KEYINPUT93), .B(n738), .Z(n739) );
  NAND2_X1 U809 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U810 ( .A(n742), .B(n741), .Z(n743) );
  NOR2_X1 U811 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U812 ( .A(KEYINPUT36), .B(n745), .ZN(n921) );
  NOR2_X1 U813 ( .A1(n777), .A2(n921), .ZN(n965) );
  NAND2_X1 U814 ( .A1(n779), .A2(n965), .ZN(n775) );
  XNOR2_X1 U815 ( .A(G1986), .B(KEYINPUT89), .ZN(n747) );
  XNOR2_X1 U816 ( .A(n747), .B(G290), .ZN(n1006) );
  INV_X1 U817 ( .A(n779), .ZN(n764) );
  NOR2_X1 U818 ( .A1(n1006), .A2(n764), .ZN(n765) );
  NAND2_X1 U819 ( .A1(G131), .A2(n914), .ZN(n749) );
  NAND2_X1 U820 ( .A1(G95), .A2(n906), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n753) );
  NAND2_X1 U822 ( .A1(G107), .A2(n908), .ZN(n751) );
  NAND2_X1 U823 ( .A1(G119), .A2(n909), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n897) );
  INV_X1 U826 ( .A(G1991), .ZN(n769) );
  NOR2_X1 U827 ( .A1(n897), .A2(n769), .ZN(n763) );
  NAND2_X1 U828 ( .A1(G141), .A2(n914), .ZN(n755) );
  NAND2_X1 U829 ( .A1(G129), .A2(n909), .ZN(n754) );
  NAND2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n759) );
  NAND2_X1 U831 ( .A1(G105), .A2(n906), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n756), .B(KEYINPUT95), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n757), .B(KEYINPUT38), .ZN(n758) );
  NOR2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n908), .A2(G117), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n902) );
  AND2_X1 U837 ( .A1(n902), .A2(G1996), .ZN(n762) );
  NOR2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n950) );
  NOR2_X1 U839 ( .A1(n950), .A2(n764), .ZN(n772) );
  XNOR2_X1 U840 ( .A(n767), .B(KEYINPUT110), .ZN(n782) );
  NOR2_X1 U841 ( .A1(G1996), .A2(n902), .ZN(n768) );
  XOR2_X1 U842 ( .A(KEYINPUT111), .B(n768), .Z(n945) );
  AND2_X1 U843 ( .A1(n769), .A2(n897), .ZN(n952) );
  NOR2_X1 U844 ( .A1(G1986), .A2(G290), .ZN(n770) );
  NOR2_X1 U845 ( .A1(n952), .A2(n770), .ZN(n771) );
  NOR2_X1 U846 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U847 ( .A1(n945), .A2(n773), .ZN(n774) );
  XNOR2_X1 U848 ( .A(n774), .B(KEYINPUT39), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U850 ( .A1(n777), .A2(n921), .ZN(n962) );
  NAND2_X1 U851 ( .A1(n778), .A2(n962), .ZN(n780) );
  NAND2_X1 U852 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U854 ( .A(n783), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U855 ( .A(G96), .ZN(G221) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G57), .ZN(G237) );
  INV_X1 U859 ( .A(G69), .ZN(G235) );
  INV_X1 U860 ( .A(G108), .ZN(G238) );
  INV_X1 U861 ( .A(G120), .ZN(G236) );
  NAND2_X1 U862 ( .A1(G94), .A2(G452), .ZN(n784) );
  XNOR2_X1 U863 ( .A(n784), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U864 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U865 ( .A(n785), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U866 ( .A(G223), .ZN(n852) );
  NAND2_X1 U867 ( .A1(n852), .A2(G567), .ZN(n786) );
  XNOR2_X1 U868 ( .A(n786), .B(KEYINPUT11), .ZN(n787) );
  XNOR2_X1 U869 ( .A(KEYINPUT69), .B(n787), .ZN(G234) );
  INV_X1 U870 ( .A(G860), .ZN(n795) );
  OR2_X1 U871 ( .A1(n994), .A2(n795), .ZN(G153) );
  INV_X1 U872 ( .A(G868), .ZN(n792) );
  NOR2_X1 U873 ( .A1(G171), .A2(n792), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT73), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n792), .A2(n996), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(G284) );
  NOR2_X1 U877 ( .A1(G868), .A2(G299), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT76), .ZN(n794) );
  NOR2_X1 U879 ( .A1(n792), .A2(G286), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(G297) );
  NAND2_X1 U881 ( .A1(n795), .A2(G559), .ZN(n796) );
  INV_X1 U882 ( .A(n996), .ZN(n823) );
  NAND2_X1 U883 ( .A1(n796), .A2(n823), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U885 ( .A1(G868), .A2(n994), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n823), .A2(G868), .ZN(n798) );
  NOR2_X1 U887 ( .A1(G559), .A2(n798), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(G282) );
  XOR2_X1 U889 ( .A(G2100), .B(KEYINPUT78), .Z(n810) );
  NAND2_X1 U890 ( .A1(G123), .A2(n909), .ZN(n801) );
  XOR2_X1 U891 ( .A(KEYINPUT18), .B(n801), .Z(n802) );
  XNOR2_X1 U892 ( .A(n802), .B(KEYINPUT77), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G111), .A2(n908), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G135), .A2(n914), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G99), .A2(n906), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n948) );
  XNOR2_X1 U899 ( .A(G2096), .B(n948), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(G156) );
  NAND2_X1 U901 ( .A1(G93), .A2(n811), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G67), .A2(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n814), .A2(n813), .ZN(n820) );
  NAND2_X1 U904 ( .A1(G80), .A2(n815), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G55), .A2(n816), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U908 ( .A(KEYINPUT79), .B(n821), .Z(n859) );
  NOR2_X1 U909 ( .A1(G868), .A2(n859), .ZN(n822) );
  XNOR2_X1 U910 ( .A(n822), .B(KEYINPUT83), .ZN(n834) );
  NAND2_X1 U911 ( .A1(G559), .A2(n823), .ZN(n824) );
  XNOR2_X1 U912 ( .A(n994), .B(n824), .ZN(n858) );
  XNOR2_X1 U913 ( .A(G166), .B(n825), .ZN(n831) );
  XNOR2_X1 U914 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n827) );
  XNOR2_X1 U915 ( .A(G290), .B(n859), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U917 ( .A(n828), .B(G305), .Z(n829) );
  XNOR2_X1 U918 ( .A(G288), .B(n829), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n831), .B(n830), .ZN(n924) );
  XOR2_X1 U920 ( .A(n858), .B(n924), .Z(n832) );
  NAND2_X1 U921 ( .A1(G868), .A2(n832), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n834), .A2(n833), .ZN(G295) );
  NAND2_X1 U923 ( .A1(G2078), .A2(G2084), .ZN(n836) );
  XOR2_X1 U924 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n835) );
  XNOR2_X1 U925 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U926 ( .A1(G2090), .A2(n837), .ZN(n838) );
  XNOR2_X1 U927 ( .A(KEYINPUT21), .B(n838), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n839), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U929 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U930 ( .A1(G236), .A2(G238), .ZN(n841) );
  NOR2_X1 U931 ( .A1(G235), .A2(G237), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U933 ( .A(KEYINPUT86), .B(n842), .ZN(n856) );
  NAND2_X1 U934 ( .A1(n856), .A2(G567), .ZN(n843) );
  XNOR2_X1 U935 ( .A(n843), .B(KEYINPUT87), .ZN(n849) );
  NOR2_X1 U936 ( .A1(G220), .A2(G219), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT22), .B(n844), .Z(n845) );
  NOR2_X1 U938 ( .A1(G218), .A2(n845), .ZN(n846) );
  XNOR2_X1 U939 ( .A(n846), .B(KEYINPUT85), .ZN(n847) );
  OR2_X1 U940 ( .A1(G221), .A2(n847), .ZN(n857) );
  AND2_X1 U941 ( .A1(G2106), .A2(n857), .ZN(n848) );
  NOR2_X1 U942 ( .A1(n849), .A2(n848), .ZN(G319) );
  INV_X1 U943 ( .A(G319), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G483), .A2(G661), .ZN(n850) );
  NOR2_X1 U945 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U946 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n852), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G661), .A2(n853), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G188) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  NOR2_X1 U955 ( .A1(n858), .A2(G860), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(G145) );
  XOR2_X1 U957 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2072), .B(G2678), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U960 ( .A(n863), .B(G2096), .Z(n865) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2090), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U963 ( .A(G2100), .B(KEYINPUT42), .Z(n867) );
  XNOR2_X1 U964 ( .A(G2078), .B(G2084), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U967 ( .A(G1961), .B(G1976), .Z(n871) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1981), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U970 ( .A(G1966), .B(G1971), .Z(n873) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U974 ( .A(KEYINPUT113), .B(G2474), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT41), .B(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G124), .A2(n909), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n908), .A2(G112), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G136), .A2(n914), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G100), .A2(n906), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G142), .A2(n914), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G106), .A2(n906), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n890), .B(KEYINPUT45), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G118), .A2(n908), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G130), .A2(n909), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(KEYINPUT114), .B(n893), .Z(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(G162), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n899) );
  XNOR2_X1 U997 ( .A(n897), .B(KEYINPUT46), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n904) );
  XOR2_X1 U1000 ( .A(G164), .B(n902), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n905), .B(n948), .Z(n920) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G103), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT115), .B(n907), .ZN(n918) );
  NAND2_X1 U1005 ( .A1(G115), .A2(n908), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G127), .A2(n909), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(KEYINPUT47), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n913), .B(KEYINPUT116), .ZN(n916) );
  NAND2_X1 U1010 ( .A1(n914), .A2(G139), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n956) );
  XNOR2_X1 U1013 ( .A(G160), .B(n956), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n922) );
  XOR2_X1 U1015 ( .A(n922), .B(n921), .Z(n923) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n923), .ZN(G395) );
  XNOR2_X1 U1017 ( .A(G171), .B(n996), .ZN(n925) );
  XNOR2_X1 U1018 ( .A(n925), .B(n924), .ZN(n927) );
  XOR2_X1 U1019 ( .A(n994), .B(G286), .Z(n926) );
  XNOR2_X1 U1020 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n928), .ZN(G397) );
  XOR2_X1 U1022 ( .A(G2451), .B(G2430), .Z(n930) );
  XNOR2_X1 U1023 ( .A(G2438), .B(G2443), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n930), .B(n929), .ZN(n936) );
  XOR2_X1 U1025 ( .A(G2435), .B(G2454), .Z(n932) );
  XNOR2_X1 U1026 ( .A(G1348), .B(G1341), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n932), .B(n931), .ZN(n934) );
  XOR2_X1 U1028 ( .A(G2446), .B(G2427), .Z(n933) );
  XNOR2_X1 U1029 ( .A(n934), .B(n933), .ZN(n935) );
  XOR2_X1 U1030 ( .A(n936), .B(n935), .Z(n937) );
  NAND2_X1 U1031 ( .A1(G14), .A2(n937), .ZN(n943) );
  NAND2_X1 U1032 ( .A1(G319), .A2(n943), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(G227), .A2(G229), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT49), .B(n938), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(G395), .A2(G397), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(G225) );
  INV_X1 U1038 ( .A(G225), .ZN(G308) );
  INV_X1 U1039 ( .A(n943), .ZN(G401) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n967) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1043 ( .A(KEYINPUT51), .B(n946), .Z(n954) );
  XOR2_X1 U1044 ( .A(G160), .B(G2084), .Z(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n961) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n955), .ZN(n958) );
  XOR2_X1 U1051 ( .A(G2072), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT50), .B(n959), .Z(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n968) );
  OR2_X1 U1058 ( .A1(KEYINPUT55), .A2(n968), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(G29), .A2(n969), .ZN(n1051) );
  INV_X1 U1060 ( .A(KEYINPUT55), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G35), .ZN(n984) );
  XOR2_X1 U1062 ( .A(n970), .B(G32), .Z(n978) );
  XNOR2_X1 U1063 ( .A(G1991), .B(G25), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G2072), .B(G33), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(G28), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(G2067), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G26), .B(n974), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G27), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1075 ( .A(G2084), .B(G34), .Z(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT54), .B(n985), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(n989), .B(n988), .ZN(n991) );
  INV_X1 U1079 ( .A(G29), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n992), .ZN(n1049) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1020) );
  XNOR2_X1 U1083 ( .A(KEYINPUT124), .B(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n1018) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT122), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G166), .B(G1971), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT123), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1010) );
  NAND2_X1 U1090 ( .A1(n703), .A2(n1002), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G299), .B(G1956), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G301), .B(G1961), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1016) );
  XNOR2_X1 U1097 ( .A(G168), .B(G1966), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT121), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1014), .B(KEYINPUT57), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1047) );
  INV_X1 U1104 ( .A(G16), .ZN(n1045) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(G4), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G19), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G1956), .B(G20), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT125), .B(G1981), .Z(n1026) );
  XNOR2_X1 U1112 ( .A(G6), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT60), .B(n1029), .Z(n1031) );
  XNOR2_X1 U1115 ( .A(G1966), .B(G21), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1041) );
  XNOR2_X1 U1117 ( .A(G1976), .B(G23), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(G22), .B(G1971), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1034), .Z(n1036) );
  XNOR2_X1 U1121 ( .A(G1986), .B(G24), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1123 ( .A(KEYINPUT58), .B(n1037), .Z(n1039) );
  XNOR2_X1 U1124 ( .A(G1961), .B(G5), .ZN(n1038) );
  NOR2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1127 ( .A(n1042), .B(KEYINPUT127), .ZN(n1043) );
  XNOR2_X1 U1128 ( .A(KEYINPUT61), .B(n1043), .ZN(n1044) );
  NAND2_X1 U1129 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1131 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  NAND2_X1 U1132 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XOR2_X1 U1133 ( .A(KEYINPUT62), .B(n1052), .Z(G311) );
  INV_X1 U1134 ( .A(G311), .ZN(G150) );
endmodule

