//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT76), .ZN(new_n203));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n205));
  OR3_X1    g004(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT78), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n203), .A2(new_n209), .A3(new_n205), .A4(new_n206), .ZN(new_n210));
  XOR2_X1   g009(.A(G141gat), .B(G148gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT79), .B(G141gat), .Z(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n202), .B2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n212), .A2(KEYINPUT81), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(new_n202), .B2(new_n204), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n221), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n214), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(KEYINPUT22), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n236), .B2(KEYINPUT29), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n229), .A3(new_n227), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(KEYINPUT84), .ZN(new_n245));
  AND2_X1   g044(.A1(G228gat), .A2(G233gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n245), .B(new_n246), .C1(new_n239), .C2(new_n243), .ZN(new_n249));
  AOI21_X1  g048(.A(G22gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(G22gat), .A3(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n250), .B2(KEYINPUT85), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n251), .A2(KEYINPUT85), .A3(new_n252), .A4(new_n256), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G226gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(G183gat), .A3(G190gat), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n266), .B1(new_n269), .B2(new_n265), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(G183gat), .B2(G190gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n272), .A2(KEYINPUT23), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(KEYINPUT23), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  AND4_X1   g077(.A1(KEYINPUT25), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n279));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n270), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(G190gat), .B1(new_n267), .B2(KEYINPUT27), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT28), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n288), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n292), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n269), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT67), .B1(new_n291), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n290), .B(new_n287), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n269), .B1(new_n299), .B2(new_n300), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n264), .B(new_n283), .C1(new_n304), .C2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n277), .A2(new_n278), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n279), .A2(new_n282), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n307), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n240), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G8gat), .B(G36gat), .Z(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT74), .ZN(new_n319));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n315), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n283), .B1(new_n304), .B2(new_n308), .ZN(new_n323));
  OAI221_X1 g122(.A(new_n236), .B1(new_n322), .B2(new_n264), .C1(new_n323), .C2(new_n311), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT30), .B1(new_n326), .B2(KEYINPUT75), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n321), .B1(new_n317), .B2(new_n324), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT30), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(new_n336), .B2(KEYINPUT69), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(KEYINPUT69), .B2(new_n336), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n339), .A2(new_n340), .A3(G134gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G113gat), .B(G120gat), .Z(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n342), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n345), .A2(KEYINPUT70), .A3(new_n346), .A4(new_n342), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n241), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n335), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n214), .A2(new_n227), .A3(new_n344), .A4(new_n351), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT82), .B1(new_n356), .B2(KEYINPUT4), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n207), .A2(KEYINPUT78), .B1(new_n212), .B2(new_n211), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n223), .B(new_n225), .C1(new_n202), .C2(new_n204), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n210), .B1(new_n362), .B2(new_n221), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT71), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(new_n360), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT71), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT71), .B1(new_n344), .B2(new_n351), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(KEYINPUT82), .A3(new_n360), .A4(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n366), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n352), .A3(new_n241), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n363), .A4(new_n364), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n360), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n373), .A2(new_n334), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n228), .A2(new_n352), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n356), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n371), .B1(new_n378), .B2(new_n335), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT86), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n333), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n370), .A3(new_n373), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT39), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n335), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n385), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT40), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n378), .B2(new_n335), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n392), .B2(new_n335), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n260), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT38), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT37), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n321), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n328), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n317), .A2(new_n324), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT37), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n403), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n372), .A2(new_n380), .A3(new_n385), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n388), .A2(new_n410), .A3(new_n411), .A4(new_n390), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n236), .B1(new_n309), .B2(new_n316), .ZN(new_n413));
  OAI221_X1 g212(.A(new_n240), .B1(new_n322), .B2(new_n264), .C1(new_n323), .C2(new_n311), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(KEYINPUT37), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n403), .B(new_n415), .C1(new_n328), .C2(new_n405), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n386), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n416), .A2(new_n417), .A3(new_n325), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n409), .B1(new_n419), .B2(KEYINPUT87), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n412), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n402), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n304), .A2(new_n308), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n314), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n359), .A2(new_n364), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n369), .A2(new_n323), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G227gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n262), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n424), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G71gat), .B(G99gat), .Z(new_n434));
  XNOR2_X1  g233(.A(G15gat), .B(G43gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT33), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n426), .A2(new_n427), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n369), .A2(new_n323), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n432), .B(new_n436), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  INV_X1    g244(.A(new_n432), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n446), .A3(new_n429), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT34), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n448), .B(new_n440), .C1(new_n433), .C2(new_n444), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n455), .A3(new_n451), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n444), .A2(new_n433), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT73), .A3(new_n448), .A4(new_n440), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(KEYINPUT36), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n417), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT83), .B1(new_n381), .B2(new_n386), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n411), .A2(new_n410), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n381), .A2(KEYINPUT83), .A3(new_n386), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n333), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n454), .B(new_n459), .C1(new_n466), .C2(new_n260), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n258), .A2(new_n259), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n456), .B2(new_n458), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n412), .A2(new_n417), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n260), .A3(new_n468), .ZN(new_n473));
  INV_X1    g272(.A(new_n333), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n452), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n423), .A2(new_n467), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G113gat), .B(G141gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G197gat), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT11), .B(G169gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT12), .Z(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT14), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT15), .A4(new_n490), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G1gat), .B2(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G8gat), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(G8gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n498), .A2(KEYINPUT17), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n496), .A2(new_n509), .A3(new_n497), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n507), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n484), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n498), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n484), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n515), .B(KEYINPUT13), .Z(new_n520));
  NOR2_X1   g319(.A1(new_n512), .A2(new_n498), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n507), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n482), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  INV_X1    g324(.A(new_n515), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT88), .B(new_n483), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n482), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n522), .A4(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n477), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G57gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G64gat), .ZN(new_n533));
  INV_X1    g332(.A(G64gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G57gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540));
  OAI21_X1  g339(.A(KEYINPUT90), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n533), .B2(new_n535), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT89), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n547));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n540), .B(new_n547), .C1(new_n537), .C2(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n541), .A2(new_n545), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(KEYINPUT21), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT92), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n512), .B1(KEYINPUT21), .B2(new_n550), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT93), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT20), .ZN(new_n559));
  XOR2_X1   g358(.A(G127gat), .B(G155gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT94), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n557), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  INV_X1    g365(.A(G99gat), .ZN(new_n567));
  INV_X1    g366(.A(G106gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT8), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G92gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n571), .B2(new_n577), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n508), .B2(new_n510), .ZN(new_n582));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n571), .A2(new_n577), .ZN(new_n586));
  INV_X1    g385(.A(new_n578), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n585), .B1(new_n499), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n565), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT96), .B1(new_n550), .B2(new_n581), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n547), .B1(new_n539), .B2(new_n540), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n542), .A2(KEYINPUT89), .A3(new_n544), .ZN(new_n605));
  AND4_X1   g404(.A1(new_n543), .A2(new_n536), .A3(new_n544), .A4(new_n538), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n590), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n550), .A2(new_n611), .A3(new_n581), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT97), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n610), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n610), .B2(new_n613), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n609), .A2(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n621), .B2(new_n616), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n590), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n541), .A2(new_n545), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n546), .A2(new_n549), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n589), .A4(new_n588), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n633), .B2(new_n612), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n618), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n616), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n626), .B1(new_n637), .B2(new_n617), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n602), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n531), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n465), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT100), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n644), .A2(new_n474), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n651), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  INV_X1    g452(.A(G8gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n644), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n333), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n651), .B2(KEYINPUT42), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n454), .A2(new_n459), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n644), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n452), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n644), .B2(new_n665), .ZN(G1326gat));
  OR3_X1    g465(.A1(new_n644), .A2(KEYINPUT102), .A3(new_n260), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT102), .B1(new_n644), .B2(new_n260), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(new_n565), .ZN(new_n673));
  INV_X1    g472(.A(new_n639), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n601), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n531), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n485), .A3(new_n465), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n477), .A2(new_n600), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n477), .A2(KEYINPUT44), .A3(new_n600), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n530), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n675), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G29gat), .B1(new_n688), .B2(new_n645), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n680), .A2(new_n689), .ZN(G1328gat));
  INV_X1    g489(.A(new_n688), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n486), .B1(new_n691), .B2(new_n333), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n486), .A3(new_n333), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n695), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n695), .B2(KEYINPUT46), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n531), .A2(new_n702), .A3(new_n452), .A4(new_n676), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT107), .Z(new_n704));
  OAI21_X1  g503(.A(G43gat), .B1(new_n688), .B2(new_n662), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1330gat));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n469), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n260), .A2(G50gat), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n709), .A2(G50gat), .B1(new_n677), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g511(.A1(new_n602), .A2(new_n530), .A3(new_n674), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n477), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n465), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(G57gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1332gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n333), .B1(new_n718), .B2(new_n534), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n534), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n714), .B2(new_n661), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n452), .A2(new_n724), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n714), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g527(.A1(new_n714), .A2(new_n469), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g529(.A1(new_n565), .A2(new_n530), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n477), .A2(new_n600), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT51), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n477), .A2(new_n734), .A3(new_n600), .A4(new_n731), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n639), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n645), .A2(G85gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n565), .A2(new_n530), .A3(new_n674), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n683), .A2(new_n684), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT110), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n683), .A2(new_n742), .A3(new_n684), .A4(new_n739), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n465), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n738), .B1(new_n744), .B2(G85gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT111), .Z(G1336gat));
  OAI21_X1  g545(.A(G92gat), .B1(new_n740), .B2(new_n474), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n474), .A2(G92gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n639), .A3(new_n735), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n741), .A2(new_n333), .A3(new_n743), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n750), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n757), .B2(KEYINPUT52), .ZN(new_n758));
  AOI211_X1 g557(.A(KEYINPUT113), .B(new_n748), .C1(new_n754), .C2(new_n756), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n751), .B1(new_n758), .B2(new_n759), .ZN(G1337gat));
  INV_X1    g559(.A(new_n736), .ZN(new_n761));
  AOI21_X1  g560(.A(G99gat), .B1(new_n761), .B2(new_n452), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n741), .A2(new_n743), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n662), .A2(new_n567), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n260), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI21_X1  g567(.A(G106gat), .B1(new_n740), .B2(new_n260), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n469), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n772), .A2(G106gat), .B1(new_n761), .B2(new_n766), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n768), .B2(new_n773), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n627), .B1(new_n637), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n620), .A2(new_n615), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n619), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n634), .A2(KEYINPUT115), .A3(new_n779), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n775), .B1(new_n621), .B2(new_n616), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n619), .A2(new_n778), .A3(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT115), .B1(new_n634), .B2(new_n779), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n786), .A2(new_n636), .A3(new_n787), .A4(KEYINPUT54), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n776), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n783), .A2(new_n777), .A3(new_n784), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n797), .B2(new_n776), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT117), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n600), .A2(new_n628), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n791), .B(new_n627), .C1(new_n637), .C2(new_n775), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n785), .B2(new_n789), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n514), .A2(new_n515), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n507), .A2(new_n521), .A3(new_n520), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n481), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n529), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT118), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(KEYINPUT118), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n801), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n800), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n674), .A2(new_n807), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n530), .A2(new_n628), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n797), .B2(new_n802), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n800), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n816), .B2(new_n600), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n673), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n602), .A2(new_n530), .A3(new_n639), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n465), .B(new_n260), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(new_n475), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n686), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n456), .A2(new_n458), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n817), .B2(new_n673), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n469), .ZN(new_n828));
  INV_X1    g627(.A(new_n825), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(KEYINPUT119), .A3(new_n465), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n474), .A3(new_n530), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n823), .B1(new_n832), .B2(new_n822), .ZN(G1340gat));
  NOR2_X1   g632(.A1(new_n674), .A2(G120gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n474), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G120gat), .B1(new_n821), .B2(new_n674), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(G1341gat));
  NAND4_X1  g638(.A1(new_n831), .A2(new_n340), .A3(new_n474), .A4(new_n565), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n821), .B2(new_n673), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  NAND2_X1  g641(.A1(new_n474), .A2(new_n600), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT121), .Z(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G134gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n831), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n821), .B2(new_n601), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  AOI21_X1  g649(.A(new_n813), .B1(new_n792), .B2(new_n815), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n601), .B1(new_n851), .B2(KEYINPUT122), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n639), .A2(new_n529), .A3(new_n806), .ZN(new_n853));
  INV_X1    g652(.A(new_n814), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n803), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n798), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n812), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n819), .B1(new_n859), .B2(new_n673), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n260), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n860), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n827), .A2(new_n260), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n865), .B(new_n866), .C1(KEYINPUT57), .C2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n661), .A2(new_n645), .A3(new_n333), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n219), .B1(new_n870), .B2(new_n686), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n869), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n215), .A3(new_n530), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT58), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n220), .A3(new_n639), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n870), .A2(new_n674), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(KEYINPUT59), .A3(new_n220), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n827), .A2(new_n864), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n859), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT124), .B(new_n812), .C1(new_n852), .C2(new_n858), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n673), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n819), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n260), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n885), .B1(new_n891), .B2(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n639), .A3(new_n869), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n880), .B1(new_n882), .B2(new_n894), .ZN(G1345gat));
  OAI21_X1  g694(.A(G155gat), .B1(new_n870), .B2(new_n673), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n872), .A2(G155gat), .A3(new_n673), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n870), .B2(new_n601), .ZN(new_n899));
  NOR4_X1   g698(.A1(new_n844), .A2(G162gat), .A3(new_n661), .A4(new_n645), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n867), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n465), .A2(new_n474), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n828), .A2(new_n452), .A3(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n296), .A3(new_n686), .ZN(new_n905));
  INV_X1    g704(.A(new_n827), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n470), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n530), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n905), .A2(new_n910), .ZN(G1348gat));
  OAI21_X1  g710(.A(G176gat), .B1(new_n904), .B2(new_n674), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n639), .A2(new_n297), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n904), .B2(new_n673), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n565), .A2(new_n917), .A3(new_n286), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n908), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n904), .B2(new_n601), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT61), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n909), .A2(new_n268), .A3(new_n600), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n892), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n661), .A2(new_n465), .A3(new_n474), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n892), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n686), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n867), .A2(new_n530), .A3(new_n927), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n930), .A2(new_n932), .B1(new_n931), .B2(new_n933), .ZN(G1352gat));
  OAI21_X1  g733(.A(G204gat), .B1(new_n929), .B2(new_n674), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n867), .A2(new_n927), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n674), .A2(G204gat), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n936), .A2(KEYINPUT62), .A3(new_n938), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(G1353gat));
  AND2_X1   g740(.A1(new_n927), .A2(new_n565), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n867), .A2(new_n231), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n944), .B(new_n231), .C1(new_n892), .C2(new_n942), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n810), .B1(new_n794), .B2(new_n799), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n600), .B1(new_n856), .B2(new_n857), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n851), .A2(KEYINPUT122), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n673), .B1(new_n949), .B2(KEYINPUT124), .ZN(new_n950));
  INV_X1    g749(.A(new_n888), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n890), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT57), .B1(new_n952), .B2(new_n469), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n942), .B1(new_n953), .B2(new_n884), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n943), .B1(new_n945), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n958), .B(new_n943), .C1(new_n945), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1354gat));
  NOR2_X1   g759(.A1(new_n601), .A2(new_n232), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n867), .A2(new_n600), .A3(new_n927), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n930), .A2(new_n961), .B1(new_n232), .B2(new_n962), .ZN(G1355gat));
endmodule


