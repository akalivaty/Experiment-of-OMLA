

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  NOR2_X1 U320 ( .A1(n490), .A2(n527), .ZN(n407) );
  XNOR2_X1 U321 ( .A(n367), .B(n366), .ZN(n371) );
  NOR2_X1 U322 ( .A1(n462), .A2(n566), .ZN(n430) );
  XOR2_X1 U323 ( .A(n293), .B(KEYINPUT22), .Z(n288) );
  AND2_X1 U324 ( .A1(n404), .A2(n403), .ZN(n289) );
  XOR2_X1 U325 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n290) );
  XNOR2_X1 U326 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n357) );
  XNOR2_X1 U327 ( .A(n358), .B(n357), .ZN(n380) );
  INV_X1 U328 ( .A(n567), .ZN(n403) );
  XNOR2_X1 U329 ( .A(n321), .B(KEYINPUT33), .ZN(n322) );
  XNOR2_X1 U330 ( .A(n323), .B(n322), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n365), .B(n364), .ZN(n366) );
  NOR2_X1 U332 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U333 ( .A(n333), .B(n332), .ZN(n334) );
  NOR2_X1 U334 ( .A1(n487), .A2(n456), .ZN(n528) );
  XNOR2_X1 U335 ( .A(n335), .B(n334), .ZN(n453) );
  XNOR2_X1 U336 ( .A(n305), .B(n304), .ZN(n462) );
  XNOR2_X1 U337 ( .A(n486), .B(n485), .ZN(n497) );
  XNOR2_X1 U338 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U339 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(G204GAT), .B(KEYINPUT23), .Z(n292) );
  NAND2_X1 U341 ( .A1(G228GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n293) );
  XNOR2_X1 U343 ( .A(G106GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n294), .B(G148GAT), .ZN(n323) );
  XNOR2_X1 U345 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n295), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U347 ( .A(n323), .B(n311), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n288), .B(n296), .ZN(n297) );
  XOR2_X1 U349 ( .A(G22GAT), .B(G155GAT), .Z(n360) );
  XOR2_X1 U350 ( .A(n297), .B(n360), .Z(n299) );
  XNOR2_X1 U351 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U353 ( .A(G162GAT), .B(KEYINPUT76), .Z(n301) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(G218GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n385) );
  XOR2_X1 U356 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n303) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n420) );
  XOR2_X1 U359 ( .A(n385), .B(n420), .Z(n304) );
  XOR2_X1 U360 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n307) );
  NAND2_X1 U361 ( .A1(G226GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n310) );
  XOR2_X1 U363 ( .A(G64GAT), .B(G92GAT), .Z(n309) );
  XNOR2_X1 U364 ( .A(G176GAT), .B(G204GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n331) );
  XOR2_X1 U366 ( .A(n310), .B(n331), .Z(n313) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(n311), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .Z(n394) );
  XOR2_X1 U370 ( .A(n314), .B(n394), .Z(n320) );
  XOR2_X1 U371 ( .A(G169GAT), .B(G8GAT), .Z(n340) );
  XNOR2_X1 U372 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n315), .B(G183GAT), .ZN(n316) );
  XOR2_X1 U374 ( .A(n316), .B(KEYINPUT18), .Z(n318) );
  XNOR2_X1 U375 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n432) );
  XNOR2_X1 U377 ( .A(n340), .B(n432), .ZN(n319) );
  XOR2_X1 U378 ( .A(n320), .B(n319), .Z(n518) );
  INV_X1 U379 ( .A(n518), .ZN(n490) );
  AND2_X1 U380 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XOR2_X1 U381 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n325) );
  XNOR2_X1 U382 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U384 ( .A(n327), .B(n326), .Z(n335) );
  XOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .Z(n393) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(n393), .ZN(n328) );
  XOR2_X1 U387 ( .A(n328), .B(KEYINPUT74), .Z(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n330) );
  XNOR2_X1 U389 ( .A(G71GAT), .B(G57GAT), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n363) );
  XNOR2_X1 U391 ( .A(n331), .B(n363), .ZN(n332) );
  INV_X1 U392 ( .A(n453), .ZN(n336) );
  XOR2_X1 U393 ( .A(n336), .B(KEYINPUT41), .Z(n549) );
  XOR2_X1 U394 ( .A(G141GAT), .B(G113GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(G50GAT), .B(G36GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U397 ( .A(n340), .B(n339), .Z(n342) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n356) );
  XOR2_X1 U400 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n344) );
  XNOR2_X1 U401 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n346) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G197GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U406 ( .A(n348), .B(n347), .Z(n354) );
  XOR2_X1 U407 ( .A(G29GAT), .B(G43GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n386) );
  XOR2_X1 U410 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n352) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(G1GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n386), .B(n359), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n567) );
  NAND2_X1 U416 ( .A1(n549), .A2(n567), .ZN(n358) );
  XOR2_X1 U417 ( .A(n360), .B(n359), .Z(n362) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n363), .B(KEYINPUT14), .ZN(n365) );
  INV_X1 U421 ( .A(KEYINPUT77), .ZN(n364) );
  XOR2_X1 U422 ( .A(G211GAT), .B(G78GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U426 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n373) );
  XNOR2_X1 U427 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(G64GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n454) );
  INV_X1 U434 ( .A(n454), .ZN(n574) );
  NOR2_X1 U435 ( .A1(n380), .A2(n574), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n381), .B(KEYINPUT114), .ZN(n397) );
  XOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n383) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U440 ( .A(n384), .B(KEYINPUT65), .Z(n388) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT10), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(G106GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U448 ( .A(n396), .B(n395), .Z(n555) );
  INV_X1 U449 ( .A(n555), .ZN(n539) );
  NAND2_X1 U450 ( .A1(n397), .A2(n539), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n398), .B(KEYINPUT47), .ZN(n405) );
  XOR2_X1 U452 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n400) );
  XNOR2_X1 U453 ( .A(KEYINPUT36), .B(n555), .ZN(n576) );
  NAND2_X1 U454 ( .A1(n574), .A2(n576), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U456 ( .A1(n401), .A2(n336), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n402), .B(KEYINPUT116), .ZN(n404) );
  NOR2_X1 U458 ( .A1(n405), .A2(n289), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n406), .B(KEYINPUT48), .ZN(n527) );
  XNOR2_X1 U460 ( .A(n407), .B(KEYINPUT54), .ZN(n428) );
  XOR2_X1 U461 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n409) );
  XNOR2_X1 U462 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n427) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G162GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G148GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n425) );
  XNOR2_X1 U471 ( .A(G127GAT), .B(G134GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n416), .B(KEYINPUT82), .ZN(n417) );
  XOR2_X1 U473 ( .A(n417), .B(KEYINPUT0), .Z(n419) );
  XNOR2_X1 U474 ( .A(G113GAT), .B(G120GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n431) );
  XOR2_X1 U476 ( .A(n420), .B(KEYINPUT4), .Z(n422) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n431), .B(n423), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U481 ( .A(n427), .B(n426), .Z(n546) );
  INV_X1 U482 ( .A(n546), .ZN(n487) );
  NAND2_X1 U483 ( .A1(n428), .A2(n487), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n429), .B(KEYINPUT64), .ZN(n566) );
  XNOR2_X1 U485 ( .A(n430), .B(n290), .ZN(n446) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n445) );
  XOR2_X1 U487 ( .A(KEYINPUT83), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G190GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n436) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n443) );
  XOR2_X1 U494 ( .A(G71GAT), .B(G176GAT), .Z(n440) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n492) );
  INV_X1 U500 ( .A(n492), .ZN(n529) );
  NAND2_X1 U501 ( .A1(n446), .A2(n529), .ZN(n561) );
  NOR2_X1 U502 ( .A1(n561), .A2(n454), .ZN(n449) );
  INV_X1 U503 ( .A(G183GAT), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT124), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(G1350GAT) );
  NOR2_X1 U506 ( .A1(n539), .A2(n561), .ZN(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n450) );
  NAND2_X1 U508 ( .A1(n453), .A2(n567), .ZN(n484) );
  NOR2_X1 U509 ( .A1(n555), .A2(n454), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT16), .B(n455), .ZN(n469) );
  XOR2_X1 U511 ( .A(n518), .B(KEYINPUT27), .Z(n460) );
  XNOR2_X1 U512 ( .A(KEYINPUT28), .B(n462), .ZN(n522) );
  OR2_X1 U513 ( .A1(n460), .A2(n522), .ZN(n456) );
  XNOR2_X1 U514 ( .A(KEYINPUT94), .B(n528), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n457), .A2(n492), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(KEYINPUT95), .ZN(n467) );
  NAND2_X1 U517 ( .A1(n462), .A2(n492), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT26), .ZN(n565) );
  NOR2_X1 U519 ( .A1(n565), .A2(n460), .ZN(n545) );
  NOR2_X1 U520 ( .A1(n490), .A2(n492), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NOR2_X1 U523 ( .A1(n545), .A2(n464), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n546), .A2(n465), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT96), .B(n468), .Z(n480) );
  NAND2_X1 U526 ( .A1(n469), .A2(n480), .ZN(n502) );
  NOR2_X1 U527 ( .A1(n484), .A2(n502), .ZN(n478) );
  NAND2_X1 U528 ( .A1(n478), .A2(n546), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT97), .Z(n473) );
  NAND2_X1 U532 ( .A1(n478), .A2(n518), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U535 ( .A1(n478), .A2(n529), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n477) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT98), .Z(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n478), .A2(n522), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n480), .A2(n576), .ZN(n481) );
  NOR2_X1 U543 ( .A1(n574), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n515) );
  NOR2_X1 U545 ( .A1(n515), .A2(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n497), .A2(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n490), .A2(n497), .ZN(n491) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U552 ( .A1(n497), .A2(n492), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT40), .B(n493), .ZN(n494) );
  INV_X1 U554 ( .A(n494), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  INV_X1 U556 ( .A(n522), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n497), .A2(n496), .ZN(n499) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n549), .Z(n560) );
  NOR2_X1 U563 ( .A1(n560), .A2(n567), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT105), .ZN(n514) );
  NOR2_X1 U565 ( .A1(n514), .A2(n502), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n546), .A2(n509), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n518), .A2(n509), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  XOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT107), .Z(n508) );
  NAND2_X1 U572 ( .A1(n509), .A2(n529), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT108), .Z(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n546), .A2(n523), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT110), .B(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT111), .Z(n520) );
  NAND2_X1 U584 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n529), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n527), .A2(n530), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n567), .A2(n534), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U596 ( .A(n534), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n560), .A2(n540), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n538) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n574), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT120), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n527), .A2(n547), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n567), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U615 ( .A1(n556), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n556), .A2(n574), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n561), .A2(n403), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n567), .A2(n577), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n577), .A2(n336), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

