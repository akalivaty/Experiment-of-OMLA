//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  INV_X1    g0008(.A(G264), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n202), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G116), .B2(G270), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT64), .B(G244), .Z(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G77), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n221), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n246), .A2(new_n248), .B1(G20), .B2(new_n203), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n206), .B2(new_n247), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  NAND4_X1  g0056(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G20), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n253), .A2(new_n258), .B1(G50), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(G50), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT67), .B(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n247), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G274), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT66), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n207), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n283), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n265), .B1(new_n293), .B2(G179), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n286), .B(KEYINPUT66), .ZN(new_n295));
  AOI211_X1 g0095(.A(new_n295), .B(new_n291), .C1(new_n279), .C2(new_n282), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n265), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n296), .B2(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n265), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n293), .A2(G200), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n301), .A2(new_n306), .A3(new_n302), .A4(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n298), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT71), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n281), .A2(new_n310), .A3(new_n289), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(G238), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT70), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n317), .A2(new_n207), .B1(new_n318), .B2(new_n274), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n319), .B2(new_n270), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n288), .B(new_n312), .C1(new_n320), .C2(new_n281), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n271), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n269), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n282), .B1(new_n324), .B2(new_n314), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n288), .A4(new_n312), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n328), .A2(KEYINPUT73), .A3(KEYINPUT14), .A4(G169), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n322), .C2(new_n327), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n322), .A2(new_n327), .A3(G179), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n329), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n248), .A2(G77), .B1(new_n251), .B2(G50), .ZN(new_n337));
  INV_X1    g0137(.A(G20), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G68), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n258), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n260), .A2(G68), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n263), .A2(G20), .A3(new_n217), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  AND4_X1   g0146(.A1(new_n340), .A2(new_n343), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT15), .B(G87), .Z(new_n349));
  AOI22_X1  g0149(.A1(new_n246), .A2(new_n251), .B1(new_n349), .B2(new_n248), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n338), .B2(new_n273), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n258), .ZN(new_n352));
  INV_X1    g0152(.A(new_n264), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n273), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n260), .A2(G77), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n277), .B2(new_n218), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n270), .A2(new_n208), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n282), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n212), .A2(new_n281), .A3(new_n289), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n288), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n363), .B2(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(G200), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n322), .A2(new_n327), .A3(G190), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n347), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n322), .B2(new_n327), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT72), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n370), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n347), .A4(new_n367), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n366), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n308), .A2(new_n348), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n266), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(G33), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n379), .A2(KEYINPUT76), .A3(G226), .A4(G1698), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n382));
  OAI21_X1  g0182(.A(G33), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n383), .A2(G226), .A3(G1698), .A4(new_n266), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(G223), .A3(new_n266), .A4(new_n271), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n380), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n282), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n288), .B1(new_n318), .B2(new_n290), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(G179), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n389), .B2(new_n282), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n331), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n267), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n247), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT75), .B1(new_n401), .B2(new_n377), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT7), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n383), .A2(new_n404), .A3(new_n266), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n383), .B2(new_n266), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n397), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n269), .A2(new_n403), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n399), .A2(new_n247), .A3(new_n400), .ZN(new_n412));
  AOI21_X1  g0212(.A(G20), .B1(new_n412), .B2(new_n268), .ZN(new_n413));
  OAI211_X1 g0213(.A(G68), .B(new_n411), .C1(new_n413), .C2(new_n408), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n397), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n417), .A3(new_n258), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n246), .A2(new_n264), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n260), .B2(new_n246), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n395), .A2(new_n421), .A3(KEYINPUT18), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n395), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n390), .A2(new_n392), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n394), .A2(G190), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n418), .A4(new_n420), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n420), .ZN(new_n432));
  INV_X1    g0232(.A(new_n258), .ZN(new_n433));
  INV_X1    g0233(.A(new_n397), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n383), .A2(new_n266), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n338), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n217), .B1(new_n436), .B2(KEYINPUT7), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n439), .B2(KEYINPUT16), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n440), .B2(new_n417), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(KEYINPUT17), .A3(new_n428), .A4(new_n427), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n363), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n362), .A2(new_n331), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n356), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n425), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n376), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(G20), .B1(G33), .B2(G283), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(G33), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT81), .B(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n258), .A2(new_n455), .A3(KEYINPUT83), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT83), .B1(new_n258), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT20), .B(new_n453), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n433), .B(new_n264), .C1(G1), .C2(new_n247), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n460), .A2(new_n461), .B1(G116), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n259), .B(G45), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(new_n281), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G270), .ZN(new_n469));
  INV_X1    g0269(.A(G274), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G257), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n317), .A2(new_n472), .B1(new_n209), .B2(new_n274), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT82), .B(G303), .Z(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n379), .B1(new_n269), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n469), .B(new_n471), .C1(new_n475), .C2(new_n281), .ZN(new_n476));
  INV_X1    g0276(.A(G190), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n454), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n264), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(G200), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n464), .A2(new_n478), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n463), .A2(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n258), .A2(new_n455), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n258), .A2(new_n455), .A3(KEYINPUT83), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n491), .B2(new_n453), .ZN(new_n492));
  INV_X1    g0292(.A(new_n461), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n481), .B(new_n486), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G169), .A3(new_n476), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n476), .A2(new_n445), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(KEYINPUT21), .A3(G169), .A4(new_n476), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n485), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n263), .A2(G20), .A3(new_n208), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n462), .A2(new_n208), .B1(KEYINPUT25), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G87), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n379), .A2(KEYINPUT22), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n479), .A2(new_n248), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n266), .A3(new_n268), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n338), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n509), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n507), .A2(new_n517), .A3(new_n508), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n504), .B1(new_n519), .B2(new_n258), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n271), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G294), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n521), .A2(new_n435), .B1(new_n247), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n282), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n468), .A2(G264), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n471), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G190), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n503), .A2(KEYINPUT25), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n520), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n379), .A2(new_n338), .A3(G68), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n313), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G20), .B1(new_n314), .B2(KEYINPUT19), .ZN(new_n535));
  NOR3_X1   g0335(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n532), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n258), .ZN(new_n538));
  INV_X1    g0338(.A(new_n349), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n353), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n540), .C1(new_n539), .C2(new_n462), .ZN(new_n541));
  INV_X1    g0341(.A(G250), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n470), .B1(new_n542), .B2(KEYINPUT80), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n259), .A3(G45), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT80), .B(G250), .C1(new_n284), .C2(G1), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n282), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n271), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n435), .B1(new_n247), .B2(new_n454), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n282), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n331), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n445), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(G200), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n537), .A2(new_n258), .B1(new_n353), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n463), .A2(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(G190), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n520), .A2(new_n530), .B1(new_n331), .B2(new_n526), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n527), .A2(new_n445), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n379), .A2(KEYINPUT78), .A3(G244), .A4(new_n271), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n271), .A2(G244), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n435), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT79), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT79), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n563), .A2(new_n566), .A3(new_n571), .A4(new_n567), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n275), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n569), .A2(new_n570), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n282), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n468), .A2(G257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n471), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n331), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n574), .B2(new_n282), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n445), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n264), .A2(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(KEYINPUT6), .B2(G97), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n208), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G107), .A3(new_n586), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(G20), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n251), .A2(G77), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n411), .B1(new_n413), .B2(new_n408), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n593), .C1(new_n208), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n583), .B1(new_n595), .B2(new_n258), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n452), .B2(new_n462), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n580), .A2(new_n582), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n581), .A2(G190), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n462), .A2(new_n452), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n583), .B(new_n600), .C1(new_n595), .C2(new_n258), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n601), .C1(new_n369), .C2(new_n581), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n562), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n450), .A2(new_n502), .A3(new_n531), .A4(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n448), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n372), .A2(new_n347), .A3(new_n367), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n348), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n425), .B1(new_n608), .B2(new_n443), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n305), .A2(new_n307), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n298), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n450), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n557), .B1(new_n369), .B2(new_n549), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n555), .A2(new_n615), .A3(new_n556), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n555), .B2(new_n556), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n553), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n601), .B1(new_n445), .B2(new_n581), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n580), .A4(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT26), .B1(new_n598), .B2(new_n559), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n553), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n520), .A2(new_n530), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n526), .A2(new_n331), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n561), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n618), .A2(new_n531), .A3(new_n553), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n598), .A4(new_n602), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n611), .B1(new_n612), .B2(new_n636), .ZN(G369));
  NOR2_X1   g0437(.A1(new_n262), .A2(G20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n259), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n464), .B2(new_n481), .ZN(new_n646));
  MUX2_X1   g0446(.A(new_n502), .B(new_n501), .S(new_n646), .Z(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT87), .Z(new_n648));
  INV_X1    g0448(.A(new_n628), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n645), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n626), .A2(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n531), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n628), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n648), .A2(G330), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n501), .A2(new_n645), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n649), .B2(new_n645), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT88), .Z(G399));
  INV_X1    g0460(.A(new_n222), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G1), .ZN(new_n664));
  INV_X1    g0464(.A(G116), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n536), .A2(new_n665), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n664), .A2(new_n666), .B1(new_n226), .B2(new_n663), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT29), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n598), .A2(KEYINPUT26), .A3(new_n559), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n598), .B2(new_n619), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n553), .A4(new_n631), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n672), .B2(new_n645), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n598), .A2(new_n602), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT86), .A3(new_n629), .A4(new_n630), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n631), .A2(new_n632), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n644), .B1(new_n677), .B2(new_n625), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n524), .A2(new_n525), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(new_n476), .A3(new_n445), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n581), .A2(new_n549), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n581), .A2(KEYINPUT30), .A3(new_n549), .A4(new_n681), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n550), .A2(new_n476), .A3(new_n445), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT89), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT89), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n579), .A2(new_n687), .A3(new_n526), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n682), .A2(KEYINPUT90), .A3(new_n683), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n685), .A3(new_n689), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n644), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n691), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n603), .A2(new_n502), .A3(new_n531), .A4(new_n645), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n679), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n668), .B1(new_n703), .B2(G1), .ZN(G364));
  NAND2_X1  g0504(.A1(new_n638), .A2(G45), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n663), .A2(G1), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n445), .A2(new_n369), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n338), .A2(G190), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G317), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G329), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n338), .A2(new_n477), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n369), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n270), .B1(new_n722), .B2(G303), .ZN(new_n723));
  INV_X1    g0523(.A(G311), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n445), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n709), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n719), .A2(new_n725), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n718), .B(new_n727), .C1(G322), .C2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n708), .A2(new_n719), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G326), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n338), .B1(new_n716), .B2(G190), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n522), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G283), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n709), .A2(new_n720), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n738), .B1(new_n736), .B2(new_n735), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n721), .A2(new_n505), .ZN(new_n742));
  INV_X1    g0542(.A(new_n740), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G107), .A2(new_n743), .B1(new_n731), .B2(G50), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n273), .B2(new_n726), .ZN(new_n745));
  INV_X1    g0545(.A(new_n734), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n742), .B(new_n745), .C1(G97), .C2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n269), .B1(new_n710), .B2(G68), .ZN(new_n748));
  INV_X1    g0548(.A(G58), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT91), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n728), .B(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n717), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G159), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT32), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n741), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n256), .B1(G20), .B2(new_n331), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n270), .A2(G355), .A3(new_n222), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n402), .A2(new_n405), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n661), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G45), .B2(new_n226), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n240), .A2(new_n284), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n758), .B1(G116), .B2(new_n222), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n757), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n756), .A2(new_n757), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n707), .B(new_n768), .C1(new_n647), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n648), .A2(G330), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n706), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n648), .A2(G330), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(G396));
  NOR2_X1   g0575(.A1(new_n448), .A2(new_n644), .ZN(new_n776));
  INV_X1    g0576(.A(new_n356), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n366), .B1(new_n777), .B2(new_n645), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n778), .B2(new_n448), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT96), .B1(new_n678), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n678), .A2(new_n779), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n780), .B(new_n781), .Z(new_n782));
  INV_X1    g0582(.A(new_n701), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n706), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n759), .ZN(new_n787));
  INV_X1    g0587(.A(new_n726), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n788), .A2(G159), .B1(new_n710), .B2(G150), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  INV_X1    g0590(.A(G143), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n732), .C1(new_n751), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n787), .B(new_n794), .C1(G58), .C2(new_n746), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n743), .A2(G68), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n202), .B2(new_n721), .C1(new_n797), .C2(new_n717), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n792), .B2(new_n793), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n479), .A2(new_n788), .B1(new_n731), .B2(G303), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n800), .B1(new_n208), .B2(new_n721), .C1(new_n522), .C2(new_n728), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n270), .B(new_n801), .C1(G283), .C2(new_n710), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n743), .A2(G87), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n724), .B2(new_n717), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G97), .B2(new_n746), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n795), .A2(new_n799), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n757), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n757), .A2(new_n764), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n807), .A2(new_n808), .B1(G77), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n779), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n706), .B(new_n811), .C1(new_n812), .C2(new_n764), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n786), .A2(new_n814), .ZN(G384));
  NAND2_X1  g0615(.A1(new_n410), .A2(new_n258), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n437), .A2(new_n438), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT16), .B1(new_n817), .B2(new_n397), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n420), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n395), .ZN(new_n820));
  INV_X1    g0620(.A(new_n642), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(new_n822), .A3(new_n429), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n395), .A2(new_n421), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT99), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n421), .B2(new_n821), .ZN(new_n827));
  AOI211_X1 g0627(.A(KEYINPUT99), .B(new_n642), .C1(new_n418), .C2(new_n420), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n429), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n824), .B1(new_n829), .B2(KEYINPUT37), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n431), .B(new_n442), .C1(new_n422), .C2(new_n423), .ZN(new_n831));
  INV_X1    g0631(.A(new_n822), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT101), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n830), .A2(new_n833), .A3(new_n836), .A4(KEYINPUT38), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n829), .A2(KEYINPUT37), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT99), .B1(new_n441), .B2(new_n642), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n421), .A2(new_n826), .A3(new_n821), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n825), .A2(new_n429), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n842), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n831), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n839), .A2(new_n845), .B1(new_n831), .B2(new_n847), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT100), .B1(new_n853), .B2(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n838), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n347), .A2(new_n645), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n348), .A2(new_n606), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n336), .A2(new_n371), .A3(new_n374), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT98), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n860), .A2(new_n861), .A3(new_n857), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n860), .B2(new_n857), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n779), .ZN(new_n865));
  NOR2_X1   g0665(.A1(KEYINPUT103), .A2(KEYINPUT31), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n695), .A2(new_n644), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n699), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n696), .A2(new_n866), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n856), .A2(KEYINPUT40), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n870), .A2(new_n699), .A3(new_n868), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n864), .A2(new_n779), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n830), .A2(new_n833), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n851), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n834), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n873), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n874), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n612), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n882), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G330), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n348), .A2(new_n644), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n879), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n835), .A2(new_n837), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n852), .B2(new_n854), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n887), .B(new_n890), .C1(new_n892), .C2(KEYINPUT39), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n635), .A2(new_n645), .A3(new_n779), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n776), .B(KEYINPUT97), .Z(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n879), .A3(new_n864), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n424), .A2(new_n642), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT102), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n893), .A2(new_n898), .A3(new_n902), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n886), .B(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n679), .A2(new_n612), .ZN(new_n906));
  INV_X1    g0706(.A(new_n611), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n905), .B(new_n908), .Z(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n259), .B2(new_n638), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n589), .A2(new_n591), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT35), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n225), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(G116), .C1(new_n912), .C2(new_n911), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n749), .B2(new_n217), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n226), .B1(G50), .B2(new_n217), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n262), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n915), .A3(new_n918), .ZN(G367));
  OAI211_X1 g0719(.A(new_n598), .B(new_n602), .C1(new_n601), .C2(new_n645), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n598), .C2(new_n645), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n924), .A2(KEYINPUT44), .A3(new_n658), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n658), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT44), .B1(new_n924), .B2(new_n658), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(new_n658), .A3(new_n927), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n925), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(new_n654), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n655), .B(new_n656), .Z(new_n934));
  XNOR2_X1  g0734(.A(new_n772), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n702), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n662), .B(KEYINPUT41), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(G1), .B(new_n705), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n654), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n924), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n616), .A2(new_n617), .A3(new_n645), .ZN(new_n942));
  MUX2_X1   g0742(.A(new_n553), .B(new_n619), .S(new_n942), .Z(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT104), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT43), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n924), .A2(new_n657), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT42), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n628), .B1(new_n922), .B2(new_n923), .ZN(new_n951));
  INV_X1    g0751(.A(new_n598), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n951), .A2(KEYINPUT106), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT106), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n645), .A3(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n946), .B(new_n948), .C1(new_n950), .C2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n950), .A2(new_n955), .A3(new_n947), .A4(new_n944), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n941), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n956), .A2(new_n958), .A3(new_n941), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT107), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n941), .C1(new_n956), .C2(new_n958), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n939), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n760), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n767), .B1(new_n222), .B2(new_n539), .C1(new_n236), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n740), .A2(new_n273), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n269), .B(new_n967), .C1(G159), .C2(new_n710), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n729), .A2(G150), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n726), .A2(new_n202), .B1(new_n717), .B2(new_n790), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G143), .B2(new_n731), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n734), .A2(new_n217), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G58), .B2(new_n722), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n726), .A2(new_n739), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n743), .A2(G97), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n711), .B2(new_n717), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(G107), .C2(new_n746), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n731), .A2(G311), .ZN(new_n979));
  INV_X1    g0779(.A(new_n751), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n474), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n787), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n722), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  INV_X1    g0783(.A(new_n710), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n721), .A2(new_n454), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n983), .B1(new_n984), .B2(new_n522), .C1(KEYINPUT46), .C2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT109), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n974), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n706), .B1(new_n989), .B2(new_n757), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n966), .B(new_n990), .C1(new_n945), .C2(new_n769), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT110), .B1(new_n964), .B2(new_n991), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(G387));
  OAI21_X1  g0796(.A(new_n760), .B1(new_n232), .B2(new_n284), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n270), .A2(new_n666), .A3(new_n222), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n217), .A2(new_n273), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n246), .A2(new_n202), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n666), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n284), .C1(KEYINPUT50), .C2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(G107), .B2(new_n222), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n655), .A2(new_n766), .B1(new_n767), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n539), .A2(new_n734), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n976), .B1(new_n202), .B2(new_n728), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(G159), .C2(new_n731), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n788), .A2(G68), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n984), .A2(new_n245), .B1(new_n717), .B2(new_n250), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G77), .B2(new_n722), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n759), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n788), .A2(new_n474), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G322), .A2(new_n731), .B1(new_n710), .B2(G311), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n751), .C2(new_n711), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT48), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n739), .B2(new_n734), .C1(new_n522), .C2(new_n721), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT111), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n759), .B1(new_n479), .B2(new_n743), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n717), .A2(new_n733), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1013), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n707), .B(new_n1006), .C1(new_n1027), .C2(new_n808), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT113), .Z(new_n1029));
  NAND2_X1  g0829(.A1(new_n935), .A2(new_n703), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n934), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n772), .B(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n702), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1033), .A3(new_n662), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n705), .A2(G1), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n935), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1029), .A2(new_n1034), .A3(new_n1036), .ZN(G393));
  INV_X1    g0837(.A(new_n933), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n663), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n933), .A2(new_n1035), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n722), .A2(G68), .B1(new_n788), .B2(new_n246), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n202), .B2(new_n984), .C1(new_n791), .C2(new_n717), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G77), .B2(new_n746), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n729), .A2(G159), .B1(new_n731), .B2(G150), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n759), .A3(new_n803), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G283), .A2(new_n722), .B1(new_n753), .B2(G322), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT115), .Z(new_n1049));
  OAI22_X1  g0849(.A1(new_n732), .A2(new_n711), .B1(new_n728), .B2(new_n724), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n710), .A2(new_n474), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n269), .B1(new_n740), .B2(new_n208), .C1(new_n522), .C2(new_n726), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n479), .B2(new_n746), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n808), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT114), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n767), .B1(new_n452), .B2(new_n222), .C1(new_n965), .C2(new_n243), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n706), .B(new_n1056), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n1057), .B2(new_n1059), .C1(new_n924), .C2(new_n769), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1040), .A2(new_n1041), .A3(new_n1061), .ZN(G390));
  NAND2_X1  g0862(.A1(new_n779), .A2(G330), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n698), .B2(new_n699), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n864), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n672), .A2(new_n645), .A3(new_n779), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n864), .B1(new_n1067), .B2(new_n895), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n887), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1069), .A3(new_n856), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n887), .B1(new_n897), .B2(new_n864), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n889), .B1(new_n856), .B2(new_n888), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1066), .B(new_n1070), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n895), .B1(new_n678), .B2(new_n779), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n864), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n890), .B1(new_n892), .B2(KEYINPUT39), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n892), .A2(new_n887), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1076), .A2(new_n1077), .B1(new_n1078), .B2(new_n1068), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1063), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n874), .A2(new_n864), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1073), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1064), .B2(new_n864), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n897), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1075), .B1(new_n883), .B2(new_n1063), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1067), .A2(new_n895), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1065), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n884), .A2(G330), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n611), .C1(new_n679), .C2(new_n612), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n662), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  INV_X1    g0896(.A(G128), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n270), .B1(new_n726), .B2(new_n1096), .C1(new_n732), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G159), .B2(new_n746), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n743), .A2(G50), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n753), .A2(G125), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n984), .A2(new_n790), .B1(new_n797), .B2(new_n728), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT53), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n721), .B2(new_n250), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n722), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n796), .B1(new_n665), .B2(new_n728), .C1(new_n522), .C2(new_n717), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G77), .B2(new_n746), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n732), .A2(new_n739), .B1(new_n726), .B2(new_n452), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n984), .A2(new_n208), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT116), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT116), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n269), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1107), .B1(new_n1114), .B2(new_n742), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n757), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n246), .B2(new_n810), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n706), .B(new_n1117), .C1(new_n1077), .C2(new_n764), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1083), .B2(new_n1035), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1095), .B1(new_n1120), .B2(new_n1121), .ZN(G378));
  NAND3_X1  g0922(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n872), .A2(G330), .A3(new_n881), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n265), .A2(new_n821), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT120), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n308), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(KEYINPUT120), .B(new_n298), .C1(new_n305), .C2(new_n307), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n308), .A2(new_n1128), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1127), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1133), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1126), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1129), .A2(new_n1131), .A3(new_n1127), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1133), .B2(new_n1130), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1125), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(G330), .A3(new_n872), .A4(new_n881), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1123), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(KEYINPUT121), .A3(new_n901), .A4(new_n903), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1035), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1140), .A2(new_n764), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n809), .A2(new_n202), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n740), .A2(new_n749), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT118), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n452), .B2(new_n984), .C1(new_n208), .C2(new_n728), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n539), .A2(new_n726), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n280), .B1(new_n273), .B2(new_n721), .C1(new_n732), .C2(new_n665), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1154), .A2(new_n972), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1157), .B(new_n787), .C1(new_n739), .C2(new_n717), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT58), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n728), .A2(new_n1097), .B1(new_n734), .B2(new_n250), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n710), .A2(G132), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n790), .B2(new_n726), .C1(new_n721), .C2(new_n1096), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G125), .C2(new_n731), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n753), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n743), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n759), .B2(G33), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1159), .B(new_n1167), .C1(G50), .C2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT119), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n706), .B1(new_n1170), .B2(new_n757), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1150), .A2(new_n1151), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1149), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1089), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1091), .B1(new_n1083), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1148), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n663), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT122), .B1(new_n904), .B2(new_n1144), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n904), .A2(new_n1144), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT122), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1146), .A2(new_n1182), .A3(new_n901), .A4(new_n903), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1173), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G375));
  NOR2_X1   g0988(.A1(new_n721), .A2(new_n452), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n728), .A2(new_n739), .B1(new_n726), .B2(new_n208), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G294), .C2(new_n731), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1007), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n753), .A2(G303), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n270), .B(new_n967), .C1(new_n479), .C2(new_n710), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n726), .A2(new_n250), .B1(new_n734), .B2(new_n202), .ZN(new_n1196));
  INV_X1    g0996(.A(G159), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n984), .A2(new_n1096), .B1(new_n1197), .B2(new_n721), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G132), .C2(new_n731), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n980), .A2(G137), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1199), .A2(new_n759), .A3(new_n1153), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n717), .A2(new_n1097), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n757), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(G68), .B2(new_n810), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n706), .B(new_n1205), .C1(new_n1075), .C2(new_n764), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1174), .B2(new_n1035), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1091), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n937), .B1(new_n1208), .B2(new_n1174), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1209), .B2(new_n1092), .ZN(G381));
  OR2_X1    g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G390), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G381), .A2(G384), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n995), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT123), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1095), .A2(new_n1119), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n995), .A2(KEYINPUT123), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1187), .A3(new_n1218), .A4(new_n1219), .ZN(G407));
  NAND3_X1  g1020(.A1(new_n1187), .A2(new_n643), .A3(new_n1218), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  NAND3_X1  g1022(.A1(G390), .A2(new_n964), .A3(new_n991), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1211), .A2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n995), .B2(G390), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1211), .B2(new_n1224), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1223), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G390), .B1(new_n964), .B2(new_n991), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1228), .A2(new_n1230), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1091), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n662), .C1(new_n1091), .C2(new_n1089), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT60), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1207), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n786), .A3(new_n814), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G384), .B(new_n1207), .C1(new_n1238), .C2(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n643), .A2(G213), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(G2897), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT124), .Z(new_n1246));
  XNOR2_X1  g1046(.A(new_n1242), .B(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1172), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1184), .B2(new_n1035), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1175), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n937), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1217), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1187), .B2(G378), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1253), .B2(new_n1244), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1248), .B1(new_n1148), .B2(new_n1035), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n662), .B1(new_n1250), .B2(KEYINPUT57), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G378), .B(new_n1255), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1218), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1242), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1243), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT62), .B1(new_n1254), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1242), .B(new_n1244), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1235), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(KEYINPUT63), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1261), .A2(new_n1243), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1247), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1270), .B(new_n1271), .C1(new_n1274), .C2(new_n1266), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(G405));
  NOR2_X1   g1076(.A1(new_n1187), .A2(new_n1217), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1258), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT127), .B1(new_n1242), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  OAI221_X1 g1083(.A(KEYINPUT127), .B1(new_n1281), .B2(new_n1242), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1283), .A2(new_n1234), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1234), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


