

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G651), .A2(n575), .ZN(n786) );
  AND2_X1 U556 ( .A1(n1001), .A2(n749), .ZN(n520) );
  OR2_X1 U557 ( .A1(n700), .A2(n690), .ZN(n521) );
  OR2_X1 U558 ( .A1(n704), .A2(n703), .ZN(n522) );
  XNOR2_X1 U559 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n602) );
  XNOR2_X1 U560 ( .A(n603), .B(n602), .ZN(n606) );
  INV_X1 U561 ( .A(n659), .ZN(n604) );
  NAND2_X1 U562 ( .A1(n521), .A2(n1008), .ZN(n691) );
  NOR2_X1 U563 ( .A1(n736), .A2(n520), .ZN(n737) );
  XNOR2_X1 U564 ( .A(n527), .B(KEYINPUT65), .ZN(n875) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n523), .ZN(n871) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n533), .Z(n785) );
  NOR2_X1 U567 ( .A1(n600), .A2(n599), .ZN(n754) );
  BUF_X1 U568 ( .A(n754), .Z(G160) );
  INV_X1 U569 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U570 ( .A1(G102), .A2(n871), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT17), .B(n524), .Z(n872) );
  NAND2_X1 U573 ( .A1(G138), .A2(n872), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n523), .A2(G2105), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G126), .A2(n875), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U578 ( .A(n528), .B(KEYINPUT67), .ZN(n876) );
  NAND2_X1 U579 ( .A1(G114), .A2(n876), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(G164) );
  INV_X1 U582 ( .A(G651), .ZN(n535) );
  NOR2_X1 U583 ( .A1(G543), .A2(n535), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n785), .A2(G65), .ZN(n538) );
  XOR2_X1 U585 ( .A(G543), .B(KEYINPUT0), .Z(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT69), .B(n534), .Z(n575) );
  OR2_X1 U587 ( .A1(n535), .A2(n575), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(n536), .Z(n782) );
  NAND2_X1 U589 ( .A1(G78), .A2(n782), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n781) );
  NAND2_X1 U592 ( .A1(n781), .A2(G91), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT72), .B(n539), .Z(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n786), .A2(G53), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G299) );
  NAND2_X1 U597 ( .A1(G64), .A2(n785), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G52), .A2(n786), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n781), .A2(G90), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT71), .B(n546), .Z(n548) );
  NAND2_X1 U602 ( .A1(G77), .A2(n782), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U606 ( .A1(G89), .A2(n781), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT4), .B(n552), .Z(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT77), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G76), .A2(n782), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n556), .ZN(n562) );
  NAND2_X1 U612 ( .A1(G63), .A2(n785), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G51), .A2(n786), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n560) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n559) );
  XNOR2_X1 U616 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n563), .ZN(G168) );
  NAND2_X1 U619 ( .A1(G88), .A2(n781), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G50), .A2(n786), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n782), .A2(G75), .ZN(n566) );
  XOR2_X1 U623 ( .A(KEYINPUT86), .B(n566), .Z(n567) );
  NOR2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n785), .A2(G62), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(G303) );
  INV_X1 U627 ( .A(G303), .ZN(G166) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G49), .A2(n786), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U632 ( .A1(n785), .A2(n573), .ZN(n574) );
  XNOR2_X1 U633 ( .A(n574), .B(KEYINPUT84), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G87), .A2(n575), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U636 ( .A1(n782), .A2(G73), .ZN(n578) );
  XNOR2_X1 U637 ( .A(n578), .B(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U638 ( .A1(G61), .A2(n785), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G48), .A2(n786), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G86), .A2(n781), .ZN(n581) );
  XNOR2_X1 U642 ( .A(KEYINPUT85), .B(n581), .ZN(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(G305) );
  NAND2_X1 U645 ( .A1(n786), .A2(G47), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G72), .A2(n782), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G85), .A2(n781), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT68), .B(n588), .Z(n589) );
  NOR2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n785), .A2(G60), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n592), .A2(n591), .ZN(G290) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NAND2_X1 U654 ( .A1(n871), .A2(G101), .ZN(n593) );
  XOR2_X1 U655 ( .A(n593), .B(KEYINPUT23), .Z(n595) );
  NAND2_X1 U656 ( .A1(n875), .A2(G125), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U658 ( .A(n596), .B(KEYINPUT66), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G137), .A2(n872), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G113), .A2(n876), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G40), .A2(n754), .ZN(n601) );
  XNOR2_X1 U663 ( .A(KEYINPUT89), .B(n601), .ZN(n705) );
  NAND2_X1 U664 ( .A1(n707), .A2(n705), .ZN(n659) );
  NAND2_X1 U665 ( .A1(G2072), .A2(n604), .ZN(n603) );
  INV_X1 U666 ( .A(G1956), .ZN(n971) );
  NOR2_X1 U667 ( .A1(n971), .A2(n604), .ZN(n605) );
  NOR2_X1 U668 ( .A1(n606), .A2(n605), .ZN(n609) );
  INV_X1 U669 ( .A(G299), .ZN(n997) );
  NOR2_X1 U670 ( .A1(n609), .A2(n997), .ZN(n608) );
  INV_X1 U671 ( .A(KEYINPUT28), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n608), .B(n607), .ZN(n646) );
  NAND2_X1 U673 ( .A1(n609), .A2(n997), .ZN(n644) );
  XNOR2_X1 U674 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n634) );
  NOR2_X1 U675 ( .A1(G1996), .A2(n634), .ZN(n620) );
  NAND2_X1 U676 ( .A1(n781), .A2(G81), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G68), .A2(n782), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n614) );
  XOR2_X1 U680 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n613) );
  XNOR2_X1 U681 ( .A(n614), .B(n613), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n785), .A2(G56), .ZN(n615) );
  XOR2_X1 U683 ( .A(KEYINPUT14), .B(n615), .Z(n616) );
  NOR2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n786), .A2(G43), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n995) );
  NOR2_X1 U687 ( .A1(n620), .A2(n995), .ZN(n632) );
  NAND2_X1 U688 ( .A1(G92), .A2(n781), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G79), .A2(n782), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U691 ( .A1(G66), .A2(n785), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G54), .A2(n786), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n628) );
  XNOR2_X1 U695 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n1004) );
  NAND2_X1 U697 ( .A1(G1348), .A2(n659), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G2067), .A2(n604), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n640) );
  NAND2_X1 U700 ( .A1(n1004), .A2(n640), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n639) );
  INV_X1 U702 ( .A(G1341), .ZN(n996) );
  NAND2_X1 U703 ( .A1(n996), .A2(n634), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n633), .A2(n659), .ZN(n637) );
  AND2_X1 U705 ( .A1(G1996), .A2(n604), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n642) );
  NOR2_X1 U709 ( .A1(n1004), .A2(n640), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U713 ( .A(KEYINPUT29), .B(n647), .Z(n651) );
  OR2_X1 U714 ( .A1(n604), .A2(G1961), .ZN(n649) );
  XNOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .ZN(n918) );
  NAND2_X1 U716 ( .A1(n604), .A2(n918), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U718 ( .A1(G171), .A2(n655), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n673) );
  NAND2_X1 U720 ( .A1(G8), .A2(n659), .ZN(n700) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n700), .ZN(n675) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n659), .ZN(n671) );
  NOR2_X1 U723 ( .A1(n675), .A2(n671), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G8), .A2(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT30), .B(n653), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U727 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT31), .B(n658), .Z(n672) );
  NOR2_X1 U730 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U731 ( .A(KEYINPUT95), .B(n660), .ZN(n663) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n700), .ZN(n661) );
  NOR2_X1 U733 ( .A1(G166), .A2(n661), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n665) );
  AND2_X1 U735 ( .A1(n672), .A2(n665), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n673), .A2(n664), .ZN(n668) );
  INV_X1 U737 ( .A(n665), .ZN(n666) );
  OR2_X1 U738 ( .A1(n666), .A2(G286), .ZN(n667) );
  AND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(G8), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U742 ( .A1(G8), .A2(n671), .ZN(n677) );
  AND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n695) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n688), .A2(n680), .ZN(n1016) );
  NAND2_X1 U750 ( .A1(n695), .A2(n1016), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT96), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G288), .A2(G1976), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n682), .B(KEYINPUT97), .ZN(n1019) );
  INV_X1 U754 ( .A(KEYINPUT98), .ZN(n683) );
  OR2_X1 U755 ( .A1(n683), .A2(n700), .ZN(n684) );
  NOR2_X1 U756 ( .A1(n1019), .A2(n684), .ZN(n685) );
  AND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U758 ( .A1(KEYINPUT33), .A2(n687), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT98), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n689), .A2(KEYINPUT33), .ZN(n690) );
  XOR2_X1 U761 ( .A(G1981), .B(G305), .Z(n1008) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n704) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U764 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U766 ( .A1(n696), .A2(n700), .ZN(n702) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(KEYINPUT93), .ZN(n698) );
  XNOR2_X1 U769 ( .A(KEYINPUT24), .B(n698), .ZN(n699) );
  OR2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  INV_X1 U772 ( .A(n705), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n749) );
  NAND2_X1 U774 ( .A1(n871), .A2(G104), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT90), .ZN(n710) );
  NAND2_X1 U776 ( .A1(G140), .A2(n872), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(KEYINPUT34), .B(n711), .ZN(n716) );
  NAND2_X1 U779 ( .A1(G128), .A2(n875), .ZN(n713) );
  NAND2_X1 U780 ( .A1(G116), .A2(n876), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U782 ( .A(KEYINPUT35), .B(n714), .Z(n715) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U784 ( .A(KEYINPUT36), .B(n717), .ZN(n889) );
  XNOR2_X1 U785 ( .A(KEYINPUT37), .B(G2067), .ZN(n747) );
  NOR2_X1 U786 ( .A1(n889), .A2(n747), .ZN(n941) );
  NAND2_X1 U787 ( .A1(n749), .A2(n941), .ZN(n745) );
  NAND2_X1 U788 ( .A1(G119), .A2(n875), .ZN(n719) );
  NAND2_X1 U789 ( .A1(G107), .A2(n876), .ZN(n718) );
  NAND2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U791 ( .A1(G95), .A2(n871), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G131), .A2(n872), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n866) );
  INV_X1 U795 ( .A(G1991), .ZN(n738) );
  NOR2_X1 U796 ( .A1(n866), .A2(n738), .ZN(n732) );
  NAND2_X1 U797 ( .A1(G129), .A2(n875), .ZN(n725) );
  NAND2_X1 U798 ( .A1(G117), .A2(n876), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U800 ( .A1(n871), .A2(G105), .ZN(n726) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(n726), .Z(n727) );
  NOR2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n872), .A2(G141), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n868) );
  AND2_X1 U805 ( .A1(n868), .A2(G1996), .ZN(n731) );
  NOR2_X1 U806 ( .A1(n732), .A2(n731), .ZN(n946) );
  XNOR2_X1 U807 ( .A(KEYINPUT91), .B(n749), .ZN(n733) );
  NOR2_X1 U808 ( .A1(n946), .A2(n733), .ZN(n742) );
  INV_X1 U809 ( .A(n742), .ZN(n734) );
  NAND2_X1 U810 ( .A1(n745), .A2(n734), .ZN(n735) );
  XNOR2_X1 U811 ( .A(n735), .B(KEYINPUT92), .ZN(n736) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n1001) );
  NAND2_X1 U813 ( .A1(n522), .A2(n737), .ZN(n752) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n868), .ZN(n956) );
  AND2_X1 U815 ( .A1(n738), .A2(n866), .ZN(n944) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n739) );
  NOR2_X1 U817 ( .A1(n944), .A2(n739), .ZN(n740) );
  XOR2_X1 U818 ( .A(KEYINPUT99), .B(n740), .Z(n741) );
  NOR2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n956), .A2(n743), .ZN(n744) );
  XNOR2_X1 U821 ( .A(n744), .B(KEYINPUT39), .ZN(n746) );
  NAND2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n889), .A2(n747), .ZN(n940) );
  NAND2_X1 U824 ( .A1(n748), .A2(n940), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U827 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  INV_X1 U830 ( .A(G132), .ZN(G219) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  XOR2_X1 U832 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n756) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U834 ( .A(n756), .B(n755), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n820) );
  NAND2_X1 U836 ( .A1(n820), .A2(G567), .ZN(n757) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n757), .Z(G234) );
  INV_X1 U838 ( .A(G860), .ZN(n763) );
  OR2_X1 U839 ( .A1(n995), .A2(n763), .ZN(G153) );
  INV_X1 U840 ( .A(G868), .ZN(n802) );
  NOR2_X1 U841 ( .A1(n802), .A2(G171), .ZN(n758) );
  XNOR2_X1 U842 ( .A(n758), .B(KEYINPUT75), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n802), .A2(n1004), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n760), .A2(n759), .ZN(G284) );
  NOR2_X1 U845 ( .A1(G286), .A2(n802), .ZN(n762) );
  NOR2_X1 U846 ( .A1(G868), .A2(G299), .ZN(n761) );
  NOR2_X1 U847 ( .A1(n762), .A2(n761), .ZN(G297) );
  NAND2_X1 U848 ( .A1(n763), .A2(G559), .ZN(n764) );
  INV_X1 U849 ( .A(n1004), .ZN(n791) );
  NAND2_X1 U850 ( .A1(n764), .A2(n791), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G559), .A2(n802), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n766), .A2(n791), .ZN(n767) );
  XNOR2_X1 U854 ( .A(n767), .B(KEYINPUT79), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n995), .A2(G868), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G282) );
  XOR2_X1 U857 ( .A(G2100), .B(KEYINPUT82), .Z(n780) );
  XOR2_X1 U858 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n771) );
  NAND2_X1 U859 ( .A1(G123), .A2(n875), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n771), .B(n770), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G99), .A2(n871), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G111), .A2(n876), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT81), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G135), .A2(n872), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n948) );
  XNOR2_X1 U868 ( .A(G2096), .B(n948), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(G156) );
  NAND2_X1 U870 ( .A1(G93), .A2(n781), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G80), .A2(n782), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G67), .A2(n785), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G55), .A2(n786), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  OR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n803) );
  NAND2_X1 U877 ( .A1(n791), .A2(G559), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(n995), .ZN(n800) );
  NOR2_X1 U879 ( .A1(G860), .A2(n800), .ZN(n793) );
  XOR2_X1 U880 ( .A(KEYINPUT83), .B(n793), .Z(n794) );
  XOR2_X1 U881 ( .A(n803), .B(n794), .Z(G145) );
  XNOR2_X1 U882 ( .A(n997), .B(KEYINPUT19), .ZN(n799) );
  XNOR2_X1 U883 ( .A(G166), .B(G305), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n795), .B(G288), .ZN(n796) );
  XOR2_X1 U885 ( .A(n803), .B(n796), .Z(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(G290), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n799), .B(n798), .ZN(n894) );
  XNOR2_X1 U888 ( .A(n800), .B(n894), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n801), .A2(G868), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n806) );
  XNOR2_X1 U893 ( .A(n806), .B(KEYINPUT87), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(KEYINPUT20), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2090), .ZN(n809) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n810), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U898 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U899 ( .A1(G483), .A2(G661), .ZN(n818) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n811) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n811), .Z(n812) );
  NOR2_X1 U902 ( .A1(G218), .A2(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G96), .A2(n813), .ZN(n914) );
  NAND2_X1 U904 ( .A1(n914), .A2(G2106), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G108), .A2(n815), .ZN(n915) );
  NAND2_X1 U908 ( .A1(n915), .A2(G567), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n826) );
  NOR2_X1 U910 ( .A1(n818), .A2(n826), .ZN(n819) );
  XNOR2_X1 U911 ( .A(n819), .B(KEYINPUT88), .ZN(n825) );
  NAND2_X1 U912 ( .A1(G36), .A2(n825), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n820), .ZN(G217) );
  INV_X1 U914 ( .A(G661), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G2), .A2(G15), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U917 ( .A(KEYINPUT104), .B(n823), .Z(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U920 ( .A(n826), .ZN(G319) );
  XOR2_X1 U921 ( .A(G2096), .B(G2100), .Z(n828) );
  XNOR2_X1 U922 ( .A(KEYINPUT42), .B(G2678), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(G2090), .Z(n830) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2072), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U927 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2084), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U930 ( .A(G1981), .B(G1956), .Z(n836) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n846) );
  XOR2_X1 U933 ( .A(KEYINPUT109), .B(G2474), .Z(n838) );
  XNOR2_X1 U934 ( .A(G1966), .B(KEYINPUT107), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n840) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1961), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n846), .B(n845), .Z(G229) );
  NAND2_X1 U943 ( .A1(G100), .A2(n871), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G136), .A2(n872), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n854) );
  NAND2_X1 U946 ( .A1(G124), .A2(n875), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n849), .B(KEYINPUT44), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT110), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G112), .A2(n876), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(G162) );
  XNOR2_X1 U952 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n872), .A2(G142), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n871), .A2(G106), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT111), .B(n855), .Z(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n863) );
  NAND2_X1 U958 ( .A1(G130), .A2(n875), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G118), .A2(n876), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n888) );
  XOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(n870) );
  XOR2_X1 U966 ( .A(G164), .B(n868), .Z(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n883) );
  NAND2_X1 U968 ( .A1(G103), .A2(n871), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G139), .A2(n872), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n882) );
  NAND2_X1 U971 ( .A1(G127), .A2(n875), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G115), .A2(n876), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT114), .B(n879), .Z(n880) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n880), .ZN(n881) );
  NOR2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n951) );
  XOR2_X1 U977 ( .A(n883), .B(n951), .Z(n885) );
  XNOR2_X1 U978 ( .A(G160), .B(G162), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U980 ( .A(n948), .B(n886), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U982 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U983 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n995), .B(G286), .ZN(n893) );
  XNOR2_X1 U985 ( .A(G171), .B(n1004), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n895) );
  XNOR2_X1 U987 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U988 ( .A1(G37), .A2(n896), .ZN(G397) );
  XNOR2_X1 U989 ( .A(KEYINPUT100), .B(G2427), .ZN(n906) );
  XOR2_X1 U990 ( .A(KEYINPUT101), .B(G2446), .Z(n898) );
  XNOR2_X1 U991 ( .A(G2435), .B(G2438), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U993 ( .A(G2454), .B(G2430), .Z(n900) );
  XNOR2_X1 U994 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2451), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(n907), .A2(G14), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(KEYINPUT102), .B(n908), .ZN(n917) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n917), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(G225) );
  XOR2_X1 U1008 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT105), .B(n916), .Z(G325) );
  XOR2_X1 U1012 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U1013 ( .A(G120), .ZN(G236) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1016 ( .A(n917), .B(KEYINPUT103), .ZN(G401) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n930) );
  XNOR2_X1 U1019 ( .A(G1991), .B(G25), .ZN(n927) );
  XNOR2_X1 U1020 ( .A(G27), .B(n918), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G1996), .B(G32), .ZN(n919) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n925), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n928), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n930), .B(n929), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT53), .B(n931), .ZN(n934) );
  XOR2_X1 U1032 ( .A(G2090), .B(KEYINPUT118), .Z(n932) );
  XNOR2_X1 U1033 ( .A(G35), .B(n932), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G34), .B(G2084), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(n935), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT55), .B(n938), .Z(n939) );
  NOR2_X1 U1039 ( .A1(G29), .A2(n939), .ZN(n968) );
  INV_X1 U1040 ( .A(n940), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G160), .B(G2084), .Z(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G2072), .B(n951), .Z(n953) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT50), .B(n954), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G2090), .B(G162), .Z(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1053 ( .A(KEYINPUT51), .B(n957), .Z(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT52), .B(n962), .ZN(n964) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(G29), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT117), .B(n966), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n1026) );
  XNOR2_X1 U1062 ( .A(G5), .B(G1961), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT125), .ZN(n983) );
  XOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .Z(n970) );
  XNOR2_X1 U1065 ( .A(G4), .B(n970), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(n996), .B(G19), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n971), .B(G20), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1071 ( .A(KEYINPUT126), .B(n976), .Z(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT60), .B(n979), .Z(n981) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G21), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n987) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n991), .ZN(n993) );
  INV_X1 U1085 ( .A(G16), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n994), .A2(G11), .ZN(n1024) );
  XOR2_X1 U1088 ( .A(G16), .B(KEYINPUT56), .Z(n1021) );
  XNOR2_X1 U1089 ( .A(n996), .B(n995), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n997), .B(G1956), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1015) );
  XOR2_X1 U1095 ( .A(n1004), .B(G1348), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(G171), .B(G1961), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT123), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1010), .B(KEYINPUT122), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT124), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
  INV_X1 U1114 ( .A(G171), .ZN(G301) );
endmodule

