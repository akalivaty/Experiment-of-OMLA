//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n207), .B(G8gat), .C1(new_n206), .C2(new_n205), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n209), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT90), .B(G8gat), .Z(new_n212));
  NAND4_X1  g011(.A1(new_n210), .A2(new_n203), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT14), .A3(new_n219), .ZN(new_n220));
  OAI221_X1 g019(.A(new_n220), .B1(KEYINPUT14), .B2(new_n219), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  AND2_X1   g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n226), .A2(KEYINPUT86), .B1(G43gat), .B2(G50gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(KEYINPUT86), .B2(new_n226), .ZN(new_n228));
  INV_X1    g027(.A(G43gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT87), .B(G50gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n224), .B1(new_n221), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n214), .B1(KEYINPUT17), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n225), .A2(new_n232), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n214), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT91), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT18), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(KEYINPUT91), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT93), .B1(new_n235), .B2(new_n214), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(new_n239), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G169gat), .B(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n246), .A3(new_n251), .A4(new_n258), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT94), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n263), .A3(new_n259), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(KEYINPUT95), .A3(new_n264), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G15gat), .B(G43gat), .Z(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  INV_X1    g077(.A(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n281), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n285), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n287), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT28), .B1(new_n287), .B2(new_n288), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n284), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n288), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n281), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n294), .A2(KEYINPUT67), .A3(G183gat), .A4(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT23), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT25), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT68), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT25), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n299), .A4(new_n297), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT64), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n288), .A3(KEYINPUT65), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n311), .A2(new_n313), .B1(new_n294), .B2(new_n296), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G169gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G176gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n299), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT25), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n291), .B1(new_n308), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT1), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n327), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n330), .B(new_n291), .C1(new_n308), .C2(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G227gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n278), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  AOI211_X1 g138(.A(KEYINPUT69), .B(new_n339), .C1(new_n332), .C2(new_n333), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n277), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n342));
  INV_X1    g141(.A(new_n333), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n322), .B1(new_n314), .B2(new_n310), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n304), .B(new_n307), .C1(new_n344), .C2(KEYINPUT25), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n330), .B1(new_n345), .B2(new_n291), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n337), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n334), .A2(new_n278), .A3(new_n337), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n276), .B(new_n341), .C1(new_n350), .C2(KEYINPUT70), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT32), .B1(new_n338), .B2(new_n340), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT73), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(new_n349), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n275), .B1(new_n358), .B2(new_n277), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT73), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n352), .B1(KEYINPUT33), .B2(new_n276), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n339), .A3(new_n333), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT34), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT74), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(G155gat), .B2(G162gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G141gat), .B(G148gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(G155gat), .B2(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n374), .C1(new_n375), .C2(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n372), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n372), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n331), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n371), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n330), .A2(new_n392), .A3(new_n383), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n330), .B2(new_n383), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n385), .A2(new_n386), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n399));
  INV_X1    g198(.A(new_n389), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n330), .A2(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT80), .B1(new_n403), .B2(new_n393), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n401), .B(new_n371), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n385), .A2(new_n386), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n408), .B2(new_n330), .ZN(new_n409));
  INV_X1    g208(.A(new_n371), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n397), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NOR2_X1   g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n416), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n421), .B2(new_n417), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G197gat), .B(G204gat), .ZN(new_n424));
  AND2_X1   g223(.A1(G211gat), .A2(G218gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(KEYINPUT22), .B2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G211gat), .B(G218gat), .Z(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT76), .ZN(new_n429));
  AND2_X1   g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n291), .C1(new_n308), .C2(new_n324), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(KEYINPUT29), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n345), .B2(new_n291), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n325), .A2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n428), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(new_n431), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT77), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n436), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n423), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n367), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n362), .A2(new_n364), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(G22gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n388), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT3), .B1(new_n428), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n408), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(G228gat), .A3(G233gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n461), .B(new_n465), .C1(new_n383), .C2(new_n462), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT31), .B(G50gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n464), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n457), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n370), .A2(new_n453), .A3(new_n455), .A4(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n454), .B1(new_n362), .B2(new_n364), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n363), .B(new_n367), .C1(new_n355), .C2(new_n361), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT6), .B1(new_n412), .B2(new_n416), .ZN(new_n481));
  INV_X1    g280(.A(new_n416), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n412), .B2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  AOI211_X1 g283(.A(new_n484), .B(new_n397), .C1(new_n407), .C2(new_n411), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n418), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR4_X1   g287(.A1(new_n488), .A2(new_n475), .A3(KEYINPUT35), .A4(new_n452), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n477), .A2(KEYINPUT35), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n478), .B2(new_n479), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n363), .B1(new_n355), .B2(new_n361), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n455), .B(KEYINPUT36), .C1(new_n494), .C2(new_n368), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n387), .A2(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT39), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n410), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n403), .A2(new_n393), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n371), .B1(new_n401), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n371), .B(new_n402), .C1(new_n408), .C2(new_n330), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT39), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n499), .B(new_n416), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT81), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n482), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n410), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(KEYINPUT40), .A3(new_n416), .A4(new_n499), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n516), .A2(new_n449), .A3(new_n450), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT83), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT37), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n436), .A2(new_n440), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n447), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT38), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT38), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n448), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n518), .B1(new_n529), .B2(new_n487), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n476), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n453), .A2(new_n475), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n496), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n270), .B1(new_n491), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(KEYINPUT8), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G99gat), .B(G106gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n233), .B2(KEYINPUT17), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n237), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n235), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n554), .A3(new_n550), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT100), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  OAI221_X1 g365(.A(new_n553), .B1(new_n560), .B2(new_n566), .C1(new_n557), .C2(new_n558), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  INV_X1    g369(.A(G71gat), .ZN(new_n571));
  INV_X1    g370(.A(G78gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(KEYINPUT96), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n576), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n214), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n580), .B(new_n582), .Z(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT97), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n568), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n544), .B(new_n576), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n544), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT102), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n595), .A2(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT101), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n610), .A3(new_n606), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n594), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n535), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n423), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g418(.A(KEYINPUT16), .B(G8gat), .Z(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n452), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(G8gat), .B1(new_n616), .B2(new_n451), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  MUX2_X1   g422(.A(new_n621), .B(new_n623), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g423(.A(G15gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n617), .A2(new_n625), .A3(new_n480), .ZN(new_n626));
  OAI21_X1  g425(.A(G15gat), .B1(new_n616), .B2(new_n496), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(G1326gat));
  NOR2_X1   g427(.A1(new_n616), .A2(new_n476), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT43), .B(G22gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1327gat));
  NOR3_X1   g430(.A1(new_n568), .A2(new_n593), .A3(new_n614), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n535), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n216), .A3(new_n423), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT45), .ZN(new_n636));
  INV_X1    g435(.A(new_n265), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n614), .A2(new_n593), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n496), .A2(KEYINPUT103), .A3(new_n533), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT103), .B1(new_n496), .B2(new_n533), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n491), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n565), .A2(KEYINPUT104), .A3(new_n567), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT104), .B1(new_n565), .B2(new_n567), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n568), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n493), .A2(new_n495), .B1(new_n531), .B2(new_n532), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n490), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT44), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n639), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G29gat), .B1(new_n654), .B2(new_n422), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n655), .ZN(G1328gat));
  NAND3_X1  g455(.A1(new_n634), .A2(new_n217), .A3(new_n452), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(KEYINPUT105), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(KEYINPUT105), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G36gat), .B1(new_n654), .B2(new_n451), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n661), .B(new_n662), .C1(new_n659), .C2(new_n657), .ZN(G1329gat));
  INV_X1    g462(.A(KEYINPUT47), .ZN(new_n664));
  INV_X1    g463(.A(new_n496), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n229), .B1(new_n653), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n480), .A2(new_n229), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n633), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT47), .B1(new_n633), .B2(new_n667), .ZN(new_n671));
  INV_X1    g470(.A(new_n639), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n534), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n650), .A2(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n677), .B2(new_n491), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n651), .A2(KEYINPUT44), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n665), .B(new_n672), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n229), .B1(new_n680), .B2(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n648), .A2(new_n652), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n665), .A4(new_n672), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n670), .B(new_n671), .C1(new_n681), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(G43gat), .A3(new_n684), .ZN(new_n687));
  INV_X1    g486(.A(new_n671), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT107), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n669), .B1(new_n685), .B2(new_n689), .ZN(G1330gat));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  INV_X1    g490(.A(new_n230), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n476), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n634), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n230), .B1(new_n653), .B2(new_n475), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n475), .B(new_n672), .C1(new_n678), .C2(new_n679), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n698), .A2(new_n696), .A3(new_n692), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n691), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701));
  INV_X1    g500(.A(new_n693), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT48), .B1(new_n633), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n230), .B1(new_n698), .B2(KEYINPUT109), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n705), .A3(new_n475), .A4(new_n672), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n701), .B(new_n703), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n692), .A3(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(new_n703), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT110), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n700), .B1(new_n707), .B2(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n614), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n594), .A2(new_n637), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n642), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n422), .B(KEYINPUT111), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n451), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n715), .B2(new_n496), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n480), .A2(new_n571), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1334gat));
  NOR2_X1   g527(.A1(new_n715), .A2(new_n476), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT113), .B(G78gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1335gat));
  INV_X1    g530(.A(new_n682), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n265), .A2(new_n592), .A3(new_n614), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n422), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n649), .A2(new_n265), .A3(new_n592), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n677), .B2(new_n491), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT51), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(new_n539), .A3(new_n423), .A4(new_n614), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(G1336gat));
  AOI21_X1  g540(.A(new_n540), .B1(new_n734), .B2(new_n452), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n738), .A2(KEYINPUT114), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n738), .A2(KEYINPUT114), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n713), .A2(G92gat), .A3(new_n451), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n744), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT52), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n747), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n753), .B2(new_n742), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n735), .B2(new_n496), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n713), .A2(G99gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n480), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1338gat));
  INV_X1    g557(.A(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n734), .B2(new_n475), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n713), .A2(new_n476), .A3(G106gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n744), .A2(new_n746), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT53), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n739), .A2(new_n761), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n767), .B2(new_n760), .ZN(G1339gat));
  NOR2_X1   g567(.A1(new_n716), .A2(new_n452), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n248), .A2(new_n250), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT116), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n240), .A2(new_n241), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n770), .B2(KEYINPUT116), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n257), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n614), .A2(new_n261), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n602), .A2(new_n776), .A3(new_n604), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n599), .B2(new_n600), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n599), .B2(new_n600), .ZN(new_n779));
  INV_X1    g578(.A(new_n610), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT55), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n613), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n784), .A3(new_n613), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n780), .A3(new_n779), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n775), .B1(new_n265), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n645), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n643), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n261), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n793), .A2(KEYINPUT117), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(KEYINPUT117), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n644), .B2(new_n645), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n593), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n594), .A2(new_n637), .A3(new_n614), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n769), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n370), .A2(new_n455), .A3(new_n476), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n637), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n792), .A2(new_n797), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n592), .ZN(new_n808));
  INV_X1    g607(.A(new_n799), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n475), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n423), .A3(new_n451), .A4(new_n480), .ZN(new_n811));
  INV_X1    g610(.A(G113gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n270), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n806), .A2(new_n813), .ZN(G1340gat));
  AOI21_X1  g613(.A(G120gat), .B1(new_n805), .B2(new_n614), .ZN(new_n815));
  INV_X1    g614(.A(G120gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n811), .A2(new_n816), .A3(new_n713), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(G1341gat));
  OAI21_X1  g617(.A(G127gat), .B1(new_n811), .B2(new_n592), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n592), .A2(G127gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n804), .B2(new_n820), .ZN(G1342gat));
  OR2_X1    g620(.A1(new_n568), .A2(G134gat), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n804), .A2(KEYINPUT56), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n811), .B2(new_n568), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT56), .B1(new_n804), .B2(new_n822), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G1343gat));
  NOR2_X1   g625(.A1(new_n665), .A2(new_n476), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n800), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G141gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n269), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n782), .B1(new_n787), .B2(new_n786), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n267), .A2(new_n268), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n649), .B1(new_n835), .B2(new_n775), .ZN(new_n836));
  INV_X1    g635(.A(new_n797), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n592), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n476), .B1(new_n838), .B2(new_n809), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n840), .B(new_n475), .C1(new_n798), .C2(new_n799), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n665), .A2(new_n422), .A3(new_n452), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n841), .A2(new_n270), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n832), .A2(G141gat), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n831), .B(new_n833), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n269), .A2(new_n830), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n800), .A2(KEYINPUT118), .A3(new_n828), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n844), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n637), .C1(new_n840), .C2(new_n839), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(G141gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n832), .B2(new_n852), .ZN(G1344gat));
  INV_X1    g652(.A(G148gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n829), .A2(new_n854), .A3(new_n614), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n796), .A2(new_n649), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n592), .B1(new_n836), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n615), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n269), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n840), .A3(new_n475), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n799), .B1(new_n807), .B2(new_n592), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n476), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n861), .A2(new_n863), .A3(new_n614), .A4(new_n843), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n856), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n856), .A2(G148gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n841), .A2(new_n844), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n614), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n855), .B1(new_n865), .B2(new_n868), .ZN(G1345gat));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  OAI21_X1  g669(.A(G155gat), .B1(new_n870), .B2(new_n592), .ZN(new_n871));
  INV_X1    g670(.A(G155gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n829), .A2(new_n872), .A3(new_n593), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n870), .B2(new_n646), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n800), .A2(G162gat), .A3(new_n568), .A4(new_n828), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n716), .A2(new_n452), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT122), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n480), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT123), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n810), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n270), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n803), .A2(new_n452), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n862), .B2(new_n423), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT120), .B(new_n422), .C1(new_n798), .C2(new_n799), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n265), .A2(G169gat), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n889), .A2(KEYINPUT121), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT121), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n884), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  AOI211_X1 g692(.A(new_n713), .B(new_n883), .C1(new_n318), .C2(new_n320), .ZN(new_n894));
  AOI21_X1  g693(.A(G176gat), .B1(new_n889), .B2(new_n614), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n882), .A2(new_n810), .A3(new_n593), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n882), .A2(new_n810), .A3(KEYINPUT124), .A4(new_n593), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G183gat), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n593), .A2(new_n287), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT60), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n901), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1350gat));
  OAI211_X1 g708(.A(new_n889), .B(new_n288), .C1(new_n644), .C2(new_n645), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n882), .A2(new_n810), .A3(new_n649), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(G190gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n288), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n912), .A2(new_n915), .B1(new_n911), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(G1351gat));
  AND2_X1   g716(.A1(new_n861), .A2(new_n863), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n880), .A2(new_n496), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G197gat), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n270), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n887), .A2(new_n888), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n827), .A2(new_n452), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT127), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n637), .A3(new_n925), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n920), .A2(new_n922), .B1(new_n921), .B2(new_n926), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n925), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n713), .A2(G204gat), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n928), .A2(KEYINPUT62), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n861), .A2(new_n863), .A3(new_n614), .A4(new_n919), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G204gat), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT62), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(G1353gat));
  OR3_X1    g733(.A1(new_n928), .A2(G211gat), .A3(new_n592), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n861), .A2(new_n863), .A3(new_n593), .A4(new_n919), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n649), .A3(new_n919), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G218gat), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n646), .A2(G218gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n928), .B2(new_n942), .ZN(G1355gat));
endmodule


