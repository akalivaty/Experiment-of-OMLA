

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n459), .B(n458), .ZN(n523) );
  XNOR2_X1 U325 ( .A(n457), .B(KEYINPUT37), .ZN(n458) );
  XNOR2_X1 U326 ( .A(n485), .B(KEYINPUT55), .ZN(n486) );
  XNOR2_X1 U327 ( .A(KEYINPUT38), .B(n461), .ZN(n508) );
  XNOR2_X1 U328 ( .A(n443), .B(n442), .ZN(n536) );
  XNOR2_X1 U329 ( .A(n404), .B(n403), .ZN(n524) );
  XOR2_X1 U330 ( .A(G155GAT), .B(KEYINPUT3), .Z(n292) );
  AND2_X1 U331 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U332 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U333 ( .A(n298), .B(n293), .ZN(n299) );
  XNOR2_X1 U334 ( .A(n396), .B(n395), .ZN(n400) );
  NOR2_X1 U335 ( .A1(n454), .A2(n453), .ZN(n494) );
  XNOR2_X1 U336 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U337 ( .A(n466), .B(KEYINPUT41), .ZN(n467) );
  AND2_X1 U338 ( .A1(n484), .A2(n483), .ZN(n574) );
  XNOR2_X1 U339 ( .A(n580), .B(n467), .ZN(n553) );
  INV_X1 U340 ( .A(G169GAT), .ZN(n487) );
  INV_X1 U341 ( .A(G29GAT), .ZN(n462) );
  XNOR2_X1 U342 ( .A(n487), .B(KEYINPUT124), .ZN(n488) );
  XNOR2_X1 U343 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U344 ( .A(n489), .B(n488), .ZN(G1348GAT) );
  XNOR2_X1 U345 ( .A(n465), .B(n464), .ZN(G1328GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n295) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G71GAT), .Z(n426) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .Z(n336) );
  XNOR2_X1 U349 ( .A(n426), .B(n336), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n300) );
  XOR2_X1 U351 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n297) );
  XNOR2_X1 U352 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n296) );
  XOR2_X1 U353 ( .A(n297), .B(n296), .Z(n298) );
  XNOR2_X1 U354 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n301), .B(KEYINPUT72), .ZN(n346) );
  XNOR2_X1 U356 ( .A(n302), .B(n346), .ZN(n308) );
  XNOR2_X1 U357 ( .A(G106GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n303), .B(G148GAT), .ZN(n418) );
  XOR2_X1 U359 ( .A(G92GAT), .B(G64GAT), .Z(n305) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT74), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U362 ( .A(G204GAT), .B(n306), .Z(n366) );
  XNOR2_X1 U363 ( .A(n418), .B(n366), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n580) );
  XOR2_X1 U365 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n310) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G29GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U368 ( .A(KEYINPUT7), .B(n311), .ZN(n332) );
  XOR2_X1 U369 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n313) );
  XNOR2_X1 U370 ( .A(KEYINPUT66), .B(KEYINPUT68), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n326) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G50GAT), .Z(n315) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(G36GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U375 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n317) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G8GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U378 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n413) );
  XOR2_X1 U380 ( .A(G113GAT), .B(G1GAT), .Z(n392) );
  XOR2_X1 U381 ( .A(n392), .B(KEYINPUT67), .Z(n321) );
  NAND2_X1 U382 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n413), .B(n322), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U387 ( .A(n332), .B(n327), .Z(n540) );
  INV_X1 U388 ( .A(n540), .ZN(n575) );
  NOR2_X1 U389 ( .A1(n580), .A2(n575), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n328), .B(KEYINPUT77), .ZN(n496) );
  XOR2_X1 U391 ( .A(KEYINPUT78), .B(KEYINPUT65), .Z(n330) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .Z(n407) );
  XOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .Z(n368) );
  XNOR2_X1 U394 ( .A(n407), .B(n368), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U396 ( .A(n331), .B(KEYINPUT11), .Z(n335) );
  INV_X1 U397 ( .A(n332), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n333), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U400 ( .A(n336), .B(G92GAT), .Z(n338) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U403 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n342) );
  XNOR2_X1 U405 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(n343), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n569) );
  XNOR2_X1 U409 ( .A(KEYINPUT36), .B(n569), .ZN(n587) );
  XOR2_X1 U410 ( .A(n346), .B(G78GAT), .Z(n348) );
  XOR2_X1 U411 ( .A(G15GAT), .B(G127GAT), .Z(n427) );
  XNOR2_X1 U412 ( .A(n427), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n353) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(G183GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n349), .B(KEYINPUT80), .ZN(n367) );
  XOR2_X1 U416 ( .A(n367), .B(KEYINPUT81), .Z(n351) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U419 ( .A(n353), .B(n352), .Z(n361) );
  XOR2_X1 U420 ( .A(G155GAT), .B(G211GAT), .Z(n355) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G1GAT), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U423 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n357) );
  XNOR2_X1 U424 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n583) );
  XNOR2_X1 U428 ( .A(G211GAT), .B(KEYINPUT92), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n362), .B(KEYINPUT21), .ZN(n363) );
  XOR2_X1 U430 ( .A(n363), .B(KEYINPUT91), .Z(n365) );
  XNOR2_X1 U431 ( .A(G197GAT), .B(G218GAT), .ZN(n364) );
  XOR2_X1 U432 ( .A(n365), .B(n364), .Z(n423) );
  XOR2_X1 U433 ( .A(n423), .B(n366), .Z(n377) );
  XOR2_X1 U434 ( .A(n368), .B(n367), .Z(n370) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U437 ( .A(n371), .B(KEYINPUT102), .Z(n375) );
  XOR2_X1 U438 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n373) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n436) );
  XNOR2_X1 U441 ( .A(n436), .B(KEYINPUT103), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n481) );
  INV_X1 U444 ( .A(KEYINPUT27), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n481), .B(n378), .ZN(n449) );
  XOR2_X1 U446 ( .A(KEYINPUT99), .B(G148GAT), .Z(n380) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(G120GAT), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U449 ( .A(G85GAT), .B(G162GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G29GAT), .B(G127GAT), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n404) );
  XOR2_X1 U453 ( .A(KEYINPUT101), .B(G57GAT), .Z(n386) );
  XNOR2_X1 U454 ( .A(KEYINPUT6), .B(KEYINPUT96), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT97), .Z(n388) );
  XNOR2_X1 U457 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n402) );
  XNOR2_X1 U460 ( .A(KEYINPUT2), .B(KEYINPUT93), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n292), .B(n391), .ZN(n406) );
  XOR2_X1 U462 ( .A(n406), .B(n392), .Z(n396) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n394) );
  INV_X1 U464 ( .A(KEYINPUT98), .ZN(n393) );
  XOR2_X1 U465 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n398) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n437) );
  XNOR2_X1 U468 ( .A(n437), .B(KEYINPUT100), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  NAND2_X1 U471 ( .A1(n449), .A2(n524), .ZN(n405) );
  XNOR2_X1 U472 ( .A(KEYINPUT104), .B(n405), .ZN(n535) );
  INV_X1 U473 ( .A(KEYINPUT28), .ZN(n425) );
  XOR2_X1 U474 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U478 ( .A(KEYINPUT89), .B(KEYINPUT95), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U480 ( .A(n412), .B(KEYINPUT23), .Z(n415) );
  XNOR2_X1 U481 ( .A(n413), .B(KEYINPUT22), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n417) );
  INV_X1 U483 ( .A(G204GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n418), .B(KEYINPUT94), .ZN(n419) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n447) );
  XNOR2_X1 U489 ( .A(n425), .B(n447), .ZN(n539) );
  XOR2_X1 U490 ( .A(G190GAT), .B(G99GAT), .Z(n429) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n441) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n431) );
  XNOR2_X1 U494 ( .A(G183GAT), .B(G176GAT), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U496 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n433) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G113GAT), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U499 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  OR2_X1 U504 ( .A1(n539), .A2(n536), .ZN(n444) );
  NOR2_X1 U505 ( .A1(n535), .A2(n444), .ZN(n454) );
  INV_X1 U506 ( .A(n481), .ZN(n526) );
  NAND2_X1 U507 ( .A1(n536), .A2(n526), .ZN(n445) );
  NAND2_X1 U508 ( .A1(n447), .A2(n445), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n446), .B(KEYINPUT25), .ZN(n451) );
  NOR2_X1 U510 ( .A1(n536), .A2(n447), .ZN(n448) );
  XNOR2_X1 U511 ( .A(KEYINPUT26), .B(n448), .ZN(n573) );
  AND2_X1 U512 ( .A1(n449), .A2(n573), .ZN(n450) );
  NOR2_X1 U513 ( .A1(n451), .A2(n450), .ZN(n452) );
  NOR2_X1 U514 ( .A1(n524), .A2(n452), .ZN(n453) );
  NOR2_X1 U515 ( .A1(n583), .A2(n494), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT108), .B(n455), .Z(n456) );
  NOR2_X1 U517 ( .A1(n587), .A2(n456), .ZN(n459) );
  INV_X1 U518 ( .A(KEYINPUT109), .ZN(n457) );
  NOR2_X1 U519 ( .A1(n496), .A2(n523), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT110), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n508), .A2(n524), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n463) );
  INV_X1 U523 ( .A(n583), .ZN(n566) );
  INV_X1 U524 ( .A(KEYINPUT64), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n553), .A2(n540), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT117), .B(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U529 ( .A1(n471), .A2(n569), .ZN(n472) );
  AND2_X1 U530 ( .A1(n566), .A2(n472), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT47), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n587), .A2(n566), .ZN(n474) );
  XOR2_X1 U533 ( .A(KEYINPUT45), .B(n474), .Z(n475) );
  NOR2_X1 U534 ( .A1(n580), .A2(n475), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n575), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n534) );
  NOR2_X1 U539 ( .A1(n481), .A2(n534), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT54), .ZN(n484) );
  INV_X1 U541 ( .A(n524), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n574), .A2(n447), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n486), .A2(n536), .ZN(n568) );
  NOR2_X1 U544 ( .A1(n575), .A2(n568), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(KEYINPUT106), .Z(n498) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n491) );
  NAND2_X1 U547 ( .A1(n583), .A2(n569), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(KEYINPUT82), .ZN(n493) );
  NOR2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U551 ( .A(KEYINPUT105), .B(n495), .ZN(n512) );
  NOR2_X1 U552 ( .A1(n496), .A2(n512), .ZN(n503) );
  NAND2_X1 U553 ( .A1(n503), .A2(n524), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n499), .Z(G1324GAT) );
  NAND2_X1 U556 ( .A1(n526), .A2(n503), .ZN(n500) );
  XNOR2_X1 U557 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U559 ( .A1(n503), .A2(n536), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n539), .A2(n503), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n504), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U563 ( .A1(n526), .A2(n508), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n508), .A2(n536), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n539), .ZN(n509) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT112), .ZN(n511) );
  XOR2_X1 U572 ( .A(KEYINPUT111), .B(n511), .Z(n514) );
  NAND2_X1 U573 ( .A1(n575), .A2(n553), .ZN(n522) );
  NOR2_X1 U574 ( .A1(n522), .A2(n512), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n519), .A2(n524), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n516) );
  NAND2_X1 U578 ( .A1(n519), .A2(n526), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n536), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U584 ( .A1(n519), .A2(n539), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n524), .A2(n529), .ZN(n525) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n529), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n529), .A2(n536), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(KEYINPUT115), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT116), .Z(n531) );
  NAND2_X1 U595 ( .A1(n529), .A2(n539), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n551) );
  NAND2_X1 U599 ( .A1(n536), .A2(n551), .ZN(n537) );
  XNOR2_X1 U600 ( .A(KEYINPUT120), .B(n537), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n540), .A2(n548), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT121), .Z(n543) );
  NAND2_X1 U605 ( .A1(n548), .A2(n553), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  NAND2_X1 U608 ( .A1(n548), .A2(n583), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  INV_X1 U612 ( .A(n569), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n551), .A2(n573), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n575), .A2(n560), .ZN(n552) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  INV_X1 U618 ( .A(n553), .ZN(n562) );
  NOR2_X1 U619 ( .A1(n562), .A2(n560), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT122), .B(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n566), .A2(n560), .ZN(n559) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n569), .A2(n560), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n568), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n568), .ZN(n567) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n579) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT59), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n586), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

