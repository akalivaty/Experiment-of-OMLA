//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT86), .B(G469), .Z(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G134), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(new_n198), .B2(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n195), .A3(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n194), .B1(new_n200), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n199), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n201), .A4(new_n203), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(G131), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(new_n209), .A3(new_n201), .A4(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n205), .A2(KEYINPUT66), .A3(G131), .A4(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT84), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G104), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n221), .A3(G104), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n227), .A2(new_n224), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n220), .A4(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n227), .A3(new_n224), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT82), .B1(new_n232), .B2(G101), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n225), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G128), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n237), .B(new_n244), .C1(new_n245), .C2(new_n241), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT10), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n231), .A2(new_n233), .ZN(new_n250));
  INV_X1    g064(.A(new_n225), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n238), .A2(G143), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n237), .A2(new_n256), .A3(new_n244), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT10), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT83), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n232), .A2(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT0), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n235), .B1(new_n262), .B2(new_n243), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT0), .B(G128), .Z(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n235), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n232), .A2(new_n266), .A3(G101), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n234), .A2(new_n270), .A3(KEYINPUT10), .A4(new_n257), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n249), .A2(new_n259), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n193), .B1(new_n219), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n234), .A2(new_n246), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n234), .A2(new_n257), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n213), .A2(new_n277), .A3(new_n214), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT12), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n215), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n247), .B1(new_n234), .B2(new_n257), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n277), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n259), .A2(new_n271), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n247), .A2(new_n248), .B1(new_n261), .B2(new_n268), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n216), .A4(new_n218), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n272), .A2(new_n280), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n193), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n285), .C2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n279), .B(new_n283), .C1(new_n219), .C2(new_n272), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n192), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n193), .A3(new_n289), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G221), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT9), .B(G234), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(new_n187), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT81), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(KEYINPUT2), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n311), .A2(new_n313), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n234), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n260), .A2(KEYINPUT4), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n231), .B2(new_n233), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n312), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n308), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G113), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT68), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n267), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n319), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n319), .B(new_n334), .C1(new_n321), .C2(new_n332), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n237), .A2(new_n256), .A3(new_n244), .A4(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n236), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n345), .A2(new_n253), .B1(new_n242), .B2(new_n243), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(KEYINPUT87), .A3(new_n341), .A4(new_n237), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n265), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT88), .B(G224), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n348), .A2(new_n355), .A3(new_n350), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n338), .A2(new_n340), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n338), .A2(new_n357), .A3(KEYINPUT89), .A4(new_n340), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n334), .B(KEYINPUT8), .ZN(new_n363));
  INV_X1    g177(.A(new_n319), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n234), .A2(new_n318), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT7), .B1(new_n355), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(new_n367), .B2(new_n355), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n348), .A2(new_n350), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n337), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n348), .A2(KEYINPUT90), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n348), .A2(KEYINPUT90), .B1(G125), .B2(new_n349), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n372), .A2(new_n373), .B1(KEYINPUT7), .B2(new_n355), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n187), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n306), .B1(new_n362), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n306), .ZN(new_n378));
  AOI211_X1 g192(.A(new_n378), .B(new_n375), .C1(new_n360), .C2(new_n361), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n305), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n304), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n382));
  NOR2_X1   g196(.A1(G237), .A2(G953), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G143), .A3(G214), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(G143), .B1(new_n383), .B2(G214), .ZN(new_n386));
  OAI21_X1  g200(.A(G131), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n209), .A3(new_n384), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n209), .B1(new_n388), .B2(new_n384), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT17), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n341), .A2(G140), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(KEYINPUT16), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT73), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n238), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT16), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(KEYINPUT73), .C1(KEYINPUT16), .C2(new_n396), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n238), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n409), .A2(KEYINPUT74), .A3(G146), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n394), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G113), .B(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(new_n223), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n396), .A2(new_n397), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(G146), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT18), .B(G131), .C1(new_n385), .C2(new_n386), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT18), .A2(G131), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n388), .A2(new_n384), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n385), .A2(new_n386), .A3(G131), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT92), .B1(new_n392), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n409), .A2(G146), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n387), .A2(new_n389), .A3(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT19), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT19), .B1(new_n396), .B2(new_n397), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n238), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n419), .ZN(new_n430));
  INV_X1    g244(.A(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n420), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT93), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n382), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(KEYINPUT20), .B(new_n435), .C1(new_n420), .C2(new_n432), .ZN(new_n438));
  INV_X1    g252(.A(G475), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n391), .A2(new_n393), .ZN(new_n440));
  INV_X1    g254(.A(new_n410), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n423), .A2(new_n403), .A3(new_n402), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n419), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n431), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n445), .B2(new_n420), .ZN(new_n446));
  OAI22_X1  g260(.A1(new_n437), .A2(new_n438), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n243), .B2(G143), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n240), .A2(KEYINPUT13), .A3(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n243), .A2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G134), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n240), .A2(G128), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n452), .A3(new_n195), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n323), .A2(G122), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n459), .A2(new_n460), .A3(new_n221), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n221), .B1(new_n459), .B2(new_n460), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G116), .B(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n221), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n456), .A2(new_n452), .A3(new_n195), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n195), .B1(new_n456), .B2(new_n452), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n459), .A2(new_n460), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n323), .A2(KEYINPUT14), .A3(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G107), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI22_X1  g287(.A1(new_n455), .A2(new_n463), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT72), .B(G217), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n352), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT94), .B1(new_n476), .B2(new_n299), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n300), .A2(new_n478), .A3(new_n352), .A4(new_n475), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n482));
  OAI221_X1 g296(.A(new_n465), .B1(new_n466), .B2(new_n467), .C1(new_n470), .C2(new_n472), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n479), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n454), .B(new_n457), .C1(new_n462), .C2(new_n461), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT95), .A4(new_n485), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n187), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G478), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n487), .A2(new_n187), .A3(new_n488), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT96), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(KEYINPUT96), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(G952), .A3(new_n352), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT21), .B(G898), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n448), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n381), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n213), .A2(new_n214), .A3(new_n265), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n195), .A2(G137), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n198), .A2(G134), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n257), .A2(new_n210), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n514), .A2(KEYINPUT30), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n330), .A2(new_n331), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT30), .B1(new_n510), .B2(new_n514), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n510), .A2(new_n517), .A3(new_n514), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n383), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT31), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n510), .A2(new_n514), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n518), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n510), .A2(KEYINPUT28), .A3(new_n517), .A4(new_n514), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n527), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n520), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n517), .B1(new_n510), .B2(new_n515), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n528), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n529), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n529), .A2(new_n537), .A3(new_n543), .A4(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT32), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n533), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n522), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n531), .A2(new_n534), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n554), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT29), .A3(new_n527), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n187), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n521), .A2(new_n555), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n536), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n535), .A2(new_n527), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT29), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G472), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n548), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n552), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G234), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n475), .B1(new_n568), .B2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n298), .A2(new_n568), .A3(G953), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n414), .A2(G146), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n409), .B2(G146), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n307), .B2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n307), .A2(G128), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n582), .A2(KEYINPUT75), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT75), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n584), .A3(new_n581), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(G110), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n243), .A2(G119), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT24), .B(G110), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n585), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n578), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n578), .A2(new_n593), .A3(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(G110), .B2(new_n587), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n441), .A2(new_n442), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n576), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT77), .ZN(new_n604));
  INV_X1    g418(.A(new_n597), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT76), .B1(new_n578), .B2(new_n593), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n601), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n598), .B2(new_n601), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n603), .B1(new_n610), .B2(new_n575), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n572), .B1(new_n611), .B2(new_n187), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT77), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n575), .B1(new_n614), .B2(new_n607), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n187), .B(new_n572), .C1(new_n615), .C2(new_n602), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n570), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n570), .A2(G902), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT79), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(KEYINPUT79), .B(new_n619), .C1(new_n615), .C2(new_n602), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n567), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT80), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n509), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n220), .ZN(G3));
  AOI21_X1  g445(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n624), .A2(new_n304), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n487), .A2(new_n638), .A3(new_n488), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n481), .A2(KEYINPUT33), .A3(new_n486), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n490), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT98), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n644), .A3(new_n640), .A4(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  INV_X1    g461(.A(new_n489), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(G478), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n489), .A2(KEYINPUT99), .A3(new_n490), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n447), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n380), .A2(new_n505), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NOR4_X1   g471(.A1(new_n380), .A2(new_n447), .A3(new_n505), .A4(new_n500), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n614), .A2(new_n607), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(KEYINPUT36), .B2(new_n576), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n610), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n619), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n618), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n602), .B1(new_n663), .B2(new_n576), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n571), .B1(new_n670), .B2(G902), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n569), .B1(new_n671), .B2(new_n616), .ZN(new_n672));
  INV_X1    g486(.A(new_n668), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT100), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n635), .A3(new_n508), .A4(new_n381), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(new_n304), .ZN(new_n679));
  INV_X1    g493(.A(new_n305), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n362), .A2(new_n376), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n378), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n362), .A2(new_n306), .A3(new_n376), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n679), .A2(new_n669), .A3(new_n674), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n567), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n502), .B1(new_n503), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n448), .A2(new_n499), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XOR2_X1   g507(.A(new_n688), .B(KEYINPUT39), .Z(new_n694));
  NAND2_X1  g508(.A1(new_n679), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n561), .A2(new_n536), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n187), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n533), .A2(new_n553), .A3(new_n522), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n527), .B1(new_n556), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n552), .A2(new_n566), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n377), .A2(new_n379), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT38), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n672), .A2(new_n673), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n433), .A2(new_n436), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT20), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n433), .A2(new_n382), .A3(new_n436), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n446), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G475), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n714), .A2(new_n716), .B1(new_n497), .B2(new_n498), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n710), .A2(new_n305), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n707), .A2(new_n709), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n698), .A2(new_n699), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NAND3_X1  g535(.A1(new_n652), .A2(new_n447), .A3(new_n689), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n652), .A2(new_n447), .A3(new_n724), .A4(new_n689), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  AOI21_X1  g543(.A(KEYINPUT32), .B1(new_n548), .B2(new_n549), .ZN(new_n730));
  INV_X1    g544(.A(new_n549), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n551), .B(new_n731), .C1(new_n546), .C2(new_n547), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n624), .B1(new_n733), .B2(new_n565), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  INV_X1    g549(.A(new_n301), .ZN(new_n736));
  INV_X1    g550(.A(new_n290), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n288), .A2(new_n279), .A3(new_n283), .A4(new_n193), .ZN(new_n738));
  AOI21_X1  g552(.A(G902), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n291), .B(new_n736), .C1(new_n739), .C2(new_n296), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n734), .A2(new_n735), .A3(new_n654), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n567), .A2(new_n654), .A3(new_n625), .A4(new_n741), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT104), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT41), .B(G113), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n745), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n734), .A2(new_n658), .A3(new_n741), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  NOR3_X1   g564(.A1(new_n380), .A2(new_n740), .A3(new_n507), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n567), .A2(new_n675), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  NAND2_X1  g567(.A1(new_n682), .A2(new_n683), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n305), .A4(new_n717), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n305), .B(new_n717), .C1(new_n377), .C2(new_n379), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n632), .A2(new_n633), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n558), .A2(new_n527), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n529), .A2(new_n543), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n731), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n740), .A2(new_n505), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n764), .A3(new_n625), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NOR3_X1   g581(.A1(new_n760), .A2(new_n710), .A3(new_n763), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n726), .A2(new_n380), .A3(new_n740), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT107), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  INV_X1    g585(.A(new_n763), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n618), .A2(new_n668), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n772), .B(new_n773), .C1(new_n633), .C2(new_n632), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n684), .A2(new_n741), .A3(new_n725), .A4(new_n723), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  INV_X1    g592(.A(new_n273), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n779), .A2(new_n289), .B1(new_n292), .B2(new_n192), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n780), .B2(G902), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n301), .B1(new_n781), .B2(new_n291), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n708), .A3(new_n305), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n567), .A2(new_n625), .A3(new_n784), .A4(new_n727), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n682), .A2(new_n305), .A3(new_n683), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n297), .A2(new_n736), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n726), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n567), .A2(new_n790), .A3(KEYINPUT42), .A4(new_n625), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n783), .A2(new_n786), .A3(new_n726), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT108), .B1(new_n734), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n787), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NAND4_X1  g611(.A1(new_n567), .A2(new_n625), .A3(new_n784), .A4(new_n691), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  OAI21_X1  g613(.A(G469), .B1(new_n780), .B2(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(KEYINPUT45), .B2(new_n780), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n296), .A2(new_n187), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n291), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n736), .B(new_n694), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT109), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n448), .A2(new_n652), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT43), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n635), .A2(new_n710), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n811));
  INV_X1    g625(.A(new_n788), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  OAI21_X1  g631(.A(new_n736), .B1(new_n804), .B2(new_n805), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT47), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n567), .A2(new_n625), .A3(new_n726), .A4(new_n788), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  INV_X1    g637(.A(new_n502), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n788), .A2(new_n740), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n734), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(KEYINPUT113), .A2(KEYINPUT48), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(G952), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n825), .A2(new_n625), .A3(new_n764), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n380), .A2(new_n740), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n830), .B(G953), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n625), .A2(new_n707), .A3(new_n502), .A4(new_n826), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n447), .A3(new_n652), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g650(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n837));
  AOI211_X1 g651(.A(new_n829), .B(new_n836), .C1(new_n827), .C2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n825), .A2(new_n768), .A3(new_n826), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n680), .A3(new_n709), .A4(new_n741), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT50), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n652), .A2(new_n447), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n839), .B(new_n841), .C1(new_n834), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n831), .A2(new_n812), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n739), .A2(new_n296), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n291), .A3(new_n302), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n819), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(KEYINPUT112), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n812), .B(new_n831), .C1(new_n820), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  OAI221_X1 g665(.A(new_n838), .B1(new_n844), .B2(new_n848), .C1(new_n851), .C2(KEYINPUT51), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT110), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n710), .A2(new_n689), .A3(new_n782), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n733), .B2(new_n705), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n853), .B1(new_n855), .B2(new_n759), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n773), .A2(new_n789), .A3(new_n688), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n853), .A2(new_n706), .A3(new_n759), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n685), .B(new_n567), .C1(new_n691), .C2(new_n727), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n777), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n706), .A2(new_n759), .A3(new_n857), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT110), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n855), .A2(new_n853), .A3(new_n759), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n777), .A4(new_n860), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n495), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n653), .B1(new_n447), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n380), .A3(new_n505), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n635), .A2(new_n873), .A3(new_n636), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n676), .A2(new_n766), .A3(new_n752), .A4(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n625), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT80), .B1(new_n567), .B2(new_n625), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n508), .B(new_n381), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n745), .A3(new_n878), .A4(new_n749), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n304), .A2(new_n447), .A3(new_n495), .A4(new_n688), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n567), .A2(new_n675), .A3(new_n880), .A4(new_n812), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n768), .A2(new_n790), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n798), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n796), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n869), .A2(new_n886), .A3(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n676), .A2(new_n766), .A3(new_n752), .A4(new_n874), .ZN(new_n889));
  INV_X1    g703(.A(new_n749), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n630), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n791), .A2(new_n792), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n794), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n883), .B1(new_n894), .B2(new_n787), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n895), .A3(new_n745), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n862), .A2(new_n868), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT111), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n887), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(KEYINPUT111), .B(new_n888), .C1(new_n896), .C2(new_n897), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n887), .A2(new_n898), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(KEYINPUT54), .B2(new_n903), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n852), .A2(new_n904), .B1(G952), .B2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n846), .A2(new_n291), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT49), .Z(new_n907));
  NOR4_X1   g721(.A1(new_n624), .A2(new_n302), .A3(new_n680), .A4(new_n808), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n707), .A3(new_n709), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(G75));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n338), .A2(new_n340), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n357), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n187), .B1(new_n887), .B2(new_n898), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT114), .B(new_n916), .C1(new_n917), .C2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT114), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n869), .B2(new_n886), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n896), .A2(new_n897), .A3(new_n888), .ZN(new_n921));
  OAI211_X1 g735(.A(G210), .B(G902), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n352), .A2(G952), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n927));
  INV_X1    g741(.A(new_n914), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n911), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n922), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n925), .B1(new_n932), .B2(new_n914), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n933), .B(KEYINPUT115), .C1(new_n923), .C2(new_n918), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G51));
  XNOR2_X1  g749(.A(new_n802), .B(KEYINPUT57), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n887), .B2(new_n898), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT116), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n737), .A2(new_n738), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(new_n936), .C1(new_n937), .C2(new_n939), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n917), .A2(new_n801), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT117), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n925), .B1(new_n945), .B2(new_n947), .ZN(G54));
  NAND3_X1  g762(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  INV_X1    g763(.A(new_n433), .ZN(new_n950));
  OR3_X1    g764(.A1(new_n949), .A2(KEYINPUT118), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT118), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n925), .B1(new_n949), .B2(new_n950), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G60));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT59), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n639), .A2(new_n640), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n937), .B2(new_n939), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(KEYINPUT119), .A3(new_n926), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n904), .A2(new_n957), .B1(new_n639), .B2(new_n640), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT119), .B1(new_n959), .B2(new_n926), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G63));
  XNOR2_X1  g777(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n965), .B(new_n966), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n887), .B2(new_n898), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n667), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n926), .B1(new_n969), .B2(new_n611), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT122), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n970), .B(new_n926), .C1(new_n611), .C2(new_n969), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n976), .A3(new_n964), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n974), .B(new_n977), .C1(new_n978), .C2(new_n975), .ZN(G66));
  NAND2_X1  g793(.A1(new_n879), .A2(new_n352), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT123), .Z(new_n981));
  INV_X1    g795(.A(new_n504), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n352), .B1(new_n982), .B2(new_n353), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n912), .B1(G898), .B2(new_n352), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(new_n538), .A2(new_n516), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n426), .A2(new_n427), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n734), .A2(new_n759), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n813), .B2(new_n814), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n861), .B1(new_n807), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n994), .A2(new_n822), .A3(new_n796), .A4(new_n798), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n352), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n352), .A2(G900), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n991), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n720), .A2(new_n777), .A3(new_n860), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n628), .A2(new_n629), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n695), .A2(new_n788), .A3(new_n872), .ZN(new_n1004));
  AOI22_X1  g818(.A1(new_n820), .A2(new_n821), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1001), .A2(new_n816), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n352), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n999), .B1(new_n1007), .B2(new_n991), .ZN(new_n1008));
  OAI21_X1  g822(.A(G953), .B1(new_n190), .B2(new_n687), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G72));
  XNOR2_X1  g824(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n633), .A2(new_n187), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n1006), .B2(new_n879), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n700), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n701), .A2(new_n562), .A3(new_n1013), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n900), .A2(new_n901), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1013), .B1(new_n995), .B2(new_n879), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n536), .A3(new_n561), .ZN(new_n1019));
  AND4_X1   g833(.A1(new_n926), .A2(new_n1015), .A3(new_n1017), .A4(new_n1019), .ZN(G57));
endmodule


