//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT74), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(G128), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n194), .B(new_n196), .C1(new_n197), .C2(KEYINPUT23), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G125), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n203), .A2(G146), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n203), .B2(new_n206), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n201), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n210), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT72), .B(G110), .Z(new_n215));
  OAI22_X1  g029(.A1(new_n198), .A2(new_n215), .B1(new_n199), .B2(new_n200), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n203), .A2(G146), .A3(new_n206), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n209), .B2(new_n218), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n192), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n192), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n219), .B2(KEYINPUT75), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n187), .B1(new_n226), .B2(G902), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  INV_X1    g042(.A(new_n187), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n225), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G234), .B2(new_n228), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT71), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n226), .A2(G902), .A3(new_n234), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n236), .A2(KEYINPUT77), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT77), .B1(new_n236), .B2(new_n238), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G140), .ZN(new_n242));
  INV_X1    g056(.A(G227), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G953), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n242), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g063(.A(G107), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G104), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(G107), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G101), .ZN(new_n254));
  AOI21_X1  g068(.A(G101), .B1(new_n247), .B2(G107), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n255), .A3(new_n251), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n195), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT0), .B(G128), .Z(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n253), .A2(new_n263), .A3(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n257), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT78), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n257), .A2(new_n267), .A3(new_n262), .A4(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n213), .A2(G143), .ZN(new_n271));
  INV_X1    g085(.A(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G146), .ZN(new_n273));
  AOI21_X1  g087(.A(G128), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(KEYINPUT1), .A3(G146), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n270), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT66), .B(new_n275), .C1(new_n258), .C2(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n258), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n248), .A2(new_n255), .A3(new_n251), .ZN(new_n284));
  INV_X1    g098(.A(G101), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n250), .A2(G104), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n252), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT79), .A3(new_n256), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n269), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n281), .B(new_n275), .C1(G128), .C2(new_n258), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n284), .A2(new_n287), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n269), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n266), .B(new_n268), .C1(new_n292), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G134), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT64), .B1(new_n298), .B2(G137), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT64), .B(new_n301), .C1(new_n298), .C2(G137), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(G137), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(new_n306), .A3(new_n302), .A4(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(KEYINPUT65), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n309), .A3(G131), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT81), .B(new_n246), .C1(new_n297), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n297), .A2(new_n311), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n281), .A2(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n295), .B1(new_n315), .B2(new_n269), .ZN(new_n316));
  INV_X1    g130(.A(new_n311), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n266), .A4(new_n268), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n246), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n293), .A2(new_n294), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n282), .B2(new_n291), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n311), .A3(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT80), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n323), .A2(new_n311), .A3(new_n326), .A4(KEYINPUT12), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n311), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n325), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n318), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n314), .A2(new_n321), .B1(new_n332), .B2(new_n245), .ZN(new_n333));
  OAI21_X1  g147(.A(G469), .B1(new_n333), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(G469), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n246), .A3(new_n318), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n246), .B1(new_n313), .B2(new_n318), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n337), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n335), .B(new_n228), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT9), .B(G234), .ZN(new_n344));
  OAI21_X1  g158(.A(G221), .B1(new_n344), .B2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G214), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n262), .A2(G125), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n277), .A2(new_n278), .B1(new_n258), .B2(new_n280), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n188), .A2(G224), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT86), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n351), .B(new_n353), .Z(new_n354));
  XOR2_X1   g168(.A(KEYINPUT2), .B(G113), .Z(new_n355));
  XNOR2_X1  g169(.A(G116), .B(G119), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n257), .A3(new_n264), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT83), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n357), .A2(new_n257), .A3(new_n360), .A4(new_n264), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n363));
  INV_X1    g177(.A(G116), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(KEYINPUT5), .A3(G119), .ZN(new_n365));
  INV_X1    g179(.A(G113), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n363), .A2(new_n367), .B1(new_n355), .B2(new_n356), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n291), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n291), .A2(new_n368), .A3(KEYINPUT84), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G122), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n362), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n362), .A2(new_n371), .A3(new_n372), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n373), .B(KEYINPUT85), .Z(new_n376));
  AOI22_X1  g190(.A1(KEYINPUT6), .A2(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n354), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT7), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n353), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n351), .B(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n373), .B(KEYINPUT8), .Z(new_n383));
  OR2_X1    g197(.A1(new_n368), .A2(new_n294), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n369), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n386), .B2(new_n374), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n389), .A3(new_n387), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n348), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n247), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT67), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G237), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G214), .A3(new_n188), .ZN(new_n403));
  AOI21_X1  g217(.A(G143), .B1(new_n403), .B2(KEYINPUT87), .ZN(new_n404));
  AOI21_X1  g218(.A(G953), .B1(new_n399), .B2(new_n401), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G214), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(KEYINPUT88), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n403), .B2(new_n272), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n407), .B2(new_n404), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n397), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n403), .A2(KEYINPUT87), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n272), .A3(new_n407), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n402), .A2(G214), .A3(new_n188), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT88), .B1(new_n416), .B2(G143), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT18), .A3(G131), .A4(new_n408), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n214), .B1(new_n213), .B2(new_n202), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n418), .A2(G131), .A3(new_n408), .ZN(new_n422));
  AOI21_X1  g236(.A(G131), .B1(new_n418), .B2(new_n408), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT17), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n418), .A2(KEYINPUT17), .A3(G131), .A4(new_n408), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  INV_X1    g240(.A(new_n208), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n217), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT89), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n396), .B(new_n421), .C1(new_n424), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n396), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n202), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n202), .B(KEYINPUT73), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n213), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n217), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n306), .B1(new_n409), .B2(new_n412), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n418), .A2(G131), .A3(new_n408), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n433), .B1(new_n434), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(G475), .A2(G902), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT20), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  INV_X1    g264(.A(new_n432), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n441), .A2(new_n442), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n425), .B(new_n430), .C1(new_n452), .C2(KEYINPUT17), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n396), .B1(new_n453), .B2(new_n421), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n228), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n448), .A2(new_n450), .B1(new_n455), .B2(G475), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n344), .A2(new_n233), .A3(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(G128), .B(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n298), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(G116), .B(G122), .Z(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(G107), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n272), .A2(G128), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(G134), .C1(KEYINPUT13), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n462), .B(new_n298), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n364), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  OAI211_X1 g287(.A(G107), .B(new_n473), .C1(new_n466), .C2(KEYINPUT14), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(new_n474), .C1(G107), .C2(new_n466), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n461), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n475), .A3(new_n461), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n460), .B1(new_n479), .B2(new_n228), .ZN(new_n480));
  INV_X1    g294(.A(new_n478), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n228), .B(new_n460), .C1(new_n481), .C2(new_n476), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n457), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n481), .A2(new_n476), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n459), .B1(new_n485), .B2(G902), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT91), .A3(new_n482), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT92), .B(G952), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G953), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(G902), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n456), .A2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n346), .A2(new_n394), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n308), .A2(new_n262), .A3(new_n310), .ZN(new_n506));
  INV_X1    g320(.A(new_n303), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n298), .A2(G137), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n307), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n282), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n506), .B2(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n357), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n357), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n405), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT31), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n515), .A2(new_n524), .A3(new_n517), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n506), .A2(new_n511), .A3(new_n516), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n516), .B1(new_n506), .B2(new_n511), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT28), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n521), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g350(.A(KEYINPUT68), .B(new_n521), .C1(new_n531), .C2(new_n533), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT69), .B1(new_n527), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n506), .A2(new_n511), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n357), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n532), .B1(new_n541), .B2(new_n517), .ZN(new_n542));
  INV_X1    g356(.A(new_n533), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT68), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n528), .A3(new_n535), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(new_n526), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n505), .B1(new_n539), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n527), .A2(new_n538), .A3(KEYINPUT69), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n545), .A2(new_n523), .A3(new_n525), .A4(new_n546), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n548), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT70), .A3(new_n505), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n515), .A2(new_n517), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n535), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n531), .A2(new_n521), .A3(new_n533), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n228), .C1(new_n561), .C2(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G472), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n503), .B1(new_n553), .B2(new_n555), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(KEYINPUT32), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n241), .B(new_n501), .C1(new_n558), .C2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  NOR3_X1   g383(.A1(new_n346), .A2(new_n240), .A3(new_n239), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n556), .A2(new_n228), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n571), .B2(G472), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n449), .B1(new_n445), .B2(new_n446), .ZN(new_n573));
  INV_X1    g387(.A(new_n446), .ZN(new_n574));
  AOI211_X1 g388(.A(KEYINPUT20), .B(new_n574), .C1(new_n432), .C2(new_n444), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n421), .B1(new_n424), .B2(new_n431), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n433), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n577), .B2(new_n432), .ZN(new_n578));
  INV_X1    g392(.A(G475), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n573), .A2(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n479), .A2(new_n458), .A3(new_n228), .ZN(new_n581));
  NAND2_X1  g395(.A1(G478), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n485), .B(KEYINPUT33), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(G478), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n498), .ZN(new_n587));
  INV_X1    g401(.A(new_n392), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n389), .B1(new_n379), .B2(new_n387), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n587), .B(new_n347), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n570), .A2(new_n572), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT34), .B(G104), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  NAND3_X1  g408(.A1(new_n448), .A2(KEYINPUT93), .A3(new_n450), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n573), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n488), .B1(new_n455), .B2(G475), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n590), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n572), .A2(new_n570), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(new_n345), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n334), .B2(new_n342), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n234), .A2(G902), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n219), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n232), .A2(new_n235), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n394), .A2(new_n500), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n572), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT37), .B(G110), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  AOI21_X1  g430(.A(KEYINPUT70), .B1(new_n556), .B2(new_n505), .ZN(new_n617));
  INV_X1    g431(.A(new_n505), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n551), .B(new_n618), .C1(new_n553), .C2(new_n555), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n556), .A2(new_n502), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(new_n504), .B1(G472), .B2(new_n564), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n611), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n494), .B1(new_n626), .B2(new_n497), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n624), .A2(new_n625), .A3(new_n393), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n595), .A2(new_n598), .A3(new_n597), .A4(new_n628), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n630), .B2(new_n394), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n623), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT95), .B(G128), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G30));
  NAND2_X1  g449(.A1(new_n621), .A2(new_n504), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n535), .B1(new_n515), .B2(new_n517), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n541), .A2(new_n517), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n228), .B1(new_n638), .B2(new_n521), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n636), .A2(new_n552), .A3(new_n557), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n588), .A2(new_n589), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n580), .A2(new_n489), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n646), .A2(new_n348), .A3(new_n610), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n627), .B(KEYINPUT39), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n605), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n642), .A2(new_n648), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT97), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G143), .ZN(G45));
  NAND3_X1  g469(.A1(new_n580), .A2(new_n585), .A3(new_n628), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n394), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n612), .B(new_n657), .C1(new_n558), .C2(new_n567), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NAND2_X1  g473(.A1(new_n313), .A2(new_n318), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n245), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT82), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n340), .A3(new_n336), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n228), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n345), .A3(new_n342), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n666), .A2(new_n586), .A3(new_n590), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n241), .B(new_n667), .C1(new_n558), .C2(new_n567), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NOR3_X1   g484(.A1(new_n666), .A2(new_n599), .A3(new_n590), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n241), .C1(new_n558), .C2(new_n567), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G116), .ZN(G18));
  NAND4_X1  g487(.A1(new_n393), .A2(new_n665), .A3(new_n345), .A4(new_n342), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n500), .A3(new_n609), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n558), .B2(new_n567), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G119), .ZN(G21));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n498), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT98), .B(G472), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n527), .A2(new_n544), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n571), .A2(new_n679), .B1(new_n502), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n236), .A2(new_n238), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT99), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n646), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n580), .A2(KEYINPUT99), .A3(new_n489), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n678), .A2(new_n681), .A3(new_n683), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  NAND2_X1  g503(.A1(new_n680), .A2(new_n502), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n553), .B2(new_n555), .ZN(new_n691));
  INV_X1    g505(.A(new_n679), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n610), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  OR3_X1    g507(.A1(new_n693), .A2(new_n656), .A3(new_n674), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  NOR3_X1   g509(.A1(new_n588), .A2(new_n589), .A3(new_n348), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n605), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT100), .B(new_n604), .C1(new_n334), .C2(new_n342), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n698), .A2(new_n656), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n636), .A2(new_n552), .A3(new_n565), .A4(new_n557), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n241), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n682), .B1(new_n622), .B2(new_n550), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n698), .A2(new_n699), .A3(new_n703), .A4(new_n656), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n702), .A2(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n306), .ZN(G33));
  NOR3_X1   g521(.A1(new_n698), .A2(new_n630), .A3(new_n699), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n701), .A3(new_n241), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G134), .ZN(G36));
  OR2_X1    g524(.A1(new_n333), .A2(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n333), .A2(KEYINPUT45), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(G469), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(G469), .A2(G902), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT46), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT102), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(KEYINPUT46), .A3(new_n714), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(new_n342), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n345), .B(new_n649), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n696), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n456), .B2(new_n585), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT103), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n580), .B(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(KEYINPUT43), .A3(new_n585), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n572), .B(new_n609), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n725), .B1(new_n730), .B2(KEYINPUT44), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n724), .B(new_n731), .C1(KEYINPUT44), .C2(new_n730), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  OAI21_X1  g547(.A(new_n345), .B1(new_n721), .B2(new_n722), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n701), .A2(new_n241), .A3(new_n656), .A4(new_n725), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G140), .ZN(G42));
  NAND3_X1  g555(.A1(new_n585), .A2(new_n347), .A3(new_n345), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n645), .A2(new_n682), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n665), .A2(new_n342), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT49), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n642), .A2(new_n743), .A3(new_n745), .A4(new_n728), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n702), .A2(new_n703), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n704), .A2(new_n705), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n668), .A2(new_n672), .A3(new_n676), .A4(new_n688), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n595), .A2(new_n597), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n486), .A2(new_n482), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT106), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(new_n628), .C1(new_n579), .C2(new_n578), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n725), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n701), .A2(new_n612), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n693), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n700), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n709), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n749), .A2(new_n750), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n568), .A2(new_n592), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n568), .A2(new_n763), .A3(new_n592), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n580), .A2(new_n753), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n590), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n570), .A2(new_n572), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n614), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n762), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT107), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n568), .A2(new_n763), .A3(new_n592), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n763), .B1(new_n568), .B2(new_n592), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n768), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n668), .A2(new_n672), .A3(new_n676), .A4(new_n688), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n706), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n759), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n612), .B1(new_n558), .B2(new_n567), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n629), .A2(new_n631), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n694), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n394), .B1(new_n685), .B2(new_n686), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n608), .A2(new_n606), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n236), .A2(new_n786), .A3(new_n628), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT108), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n609), .A2(KEYINPUT108), .A3(new_n628), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n346), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n640), .B1(new_n566), .B2(KEYINPUT32), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n785), .B(new_n791), .C1(new_n558), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n658), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n781), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n580), .A2(KEYINPUT99), .A3(new_n489), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT99), .B1(new_n580), .B2(new_n489), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n393), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n790), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n605), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n623), .A2(new_n657), .B1(new_n801), .B2(new_n641), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n693), .A2(new_n656), .A3(new_n674), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n623), .B2(new_n632), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT52), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n795), .A2(new_n805), .A3(KEYINPUT110), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n795), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n780), .A2(KEYINPUT53), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n780), .A2(new_n809), .A3(KEYINPUT111), .A4(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n802), .A2(new_n804), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT52), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n795), .A2(new_n805), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT109), .B1(new_n802), .B2(new_n804), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n780), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n812), .A2(new_n813), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT54), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n821), .B1(new_n779), .B2(new_n808), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n774), .A2(new_n759), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n774), .A2(new_n829), .A3(new_n759), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n706), .A2(new_n776), .A3(new_n821), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n819), .A2(new_n828), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n666), .A2(new_n725), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n642), .A2(new_n241), .A3(new_n494), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n727), .A2(new_n729), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n494), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n681), .A2(new_n683), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n491), .B1(new_n586), .B2(new_n837), .C1(new_n844), .C2(new_n674), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n744), .B(KEYINPUT116), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n345), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n738), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n841), .A2(new_n843), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n696), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n645), .A2(new_n347), .A3(new_n666), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT117), .Z(new_n853));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n843), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT50), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n836), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n841), .B2(new_n836), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n757), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n837), .A2(new_n580), .A3(new_n585), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n845), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n858), .A2(new_n859), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n704), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT48), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n868), .A3(new_n704), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n854), .B(KEYINPUT50), .Z(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n860), .A3(new_n862), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n847), .B1(new_n738), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n736), .A2(KEYINPUT115), .A3(new_n737), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n850), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n864), .B(new_n870), .C1(new_n877), .C2(KEYINPUT51), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n824), .B1(new_n823), .B2(KEYINPUT54), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n835), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n746), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n188), .A2(G952), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n228), .B1(new_n826), .B2(new_n832), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n377), .A2(new_n378), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n354), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT120), .Z(new_n889));
  AOI21_X1  g703(.A(new_n883), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n833), .A2(G210), .A3(G902), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT119), .B1(new_n893), .B2(new_n888), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  INV_X1    g709(.A(new_n888), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n895), .B(new_n896), .C1(new_n891), .C2(new_n892), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n890), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n900), .B(new_n890), .C1(new_n894), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(G51));
  XNOR2_X1  g716(.A(new_n833), .B(KEYINPUT54), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n714), .B(KEYINPUT57), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n663), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n713), .B(KEYINPUT122), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n884), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n883), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NAND2_X1  g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n884), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(new_n445), .ZN(new_n913));
  INV_X1    g727(.A(new_n883), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n445), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n913), .A2(new_n918), .A3(new_n914), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(G60));
  INV_X1    g734(.A(new_n584), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n582), .B(KEYINPUT59), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n903), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n914), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n835), .B2(new_n879), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n584), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n833), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n883), .B1(new_n929), .B2(new_n226), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n833), .A2(new_n608), .A3(new_n928), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT61), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n495), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n770), .A2(new_n776), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n886), .B1(G898), .B2(new_n188), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  NOR2_X1   g759(.A1(new_n513), .A2(new_n514), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n438), .Z(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n626), .B2(new_n188), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n740), .A2(new_n732), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n804), .A2(new_n658), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n749), .A2(new_n709), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n704), .A2(new_n785), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n724), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n948), .B1(new_n956), .B2(new_n188), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n654), .A2(new_n951), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n725), .B(new_n650), .C1(new_n586), .C2(new_n765), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n701), .A3(new_n241), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n949), .A2(new_n959), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n947), .B1(new_n963), .B2(new_n188), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n243), .B2(new_n626), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n942), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n955), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n517), .A3(new_n515), .A4(new_n535), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n969), .B1(new_n963), .B2(new_n970), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n637), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n974), .A3(new_n914), .ZN(new_n975));
  INV_X1    g789(.A(new_n969), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n560), .B2(new_n522), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n823), .B2(new_n977), .ZN(G57));
endmodule


