//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  XNOR2_X1  g000(.A(G183gat), .B(G211gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT97), .A2(G57gat), .A3(G64gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n206));
  INV_X1    g005(.A(G64gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT96), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT98), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n211), .B(KEYINPUT96), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT98), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT99), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G57gat), .B(G64gat), .Z(new_n221));
  AOI21_X1  g020(.A(new_n204), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(KEYINPUT98), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(new_n214), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT99), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT21), .ZN(new_n229));
  AND2_X1   g028(.A1(G231gat), .A2(G233gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G127gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n203), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n203), .A3(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT88), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G1gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT89), .ZN(new_n244));
  XNOR2_X1  g043(.A(G15gat), .B(G22gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT87), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n245), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n239), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT90), .B(G8gat), .Z(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT91), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n243), .A2(KEYINPUT89), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n243), .A2(KEYINPUT89), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n246), .A2(G1gat), .ZN(new_n257));
  OAI21_X1  g056(.A(G8gat), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n247), .A2(new_n259), .A3(new_n250), .A4(new_n251), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(KEYINPUT21), .B2(new_n228), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT100), .Z(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n264));
  INV_X1    g063(.A(G155gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n266), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n236), .A2(new_n237), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n263), .B(new_n266), .ZN(new_n270));
  INV_X1    g069(.A(new_n237), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n235), .ZN(new_n272));
  NOR2_X1   g071(.A1(G29gat), .A2(G36gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT14), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G29gat), .A2(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT86), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT15), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(KEYINPUT15), .A3(new_n277), .ZN(new_n281));
  XNOR2_X1  g080(.A(G43gat), .B(G50gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G85gat), .A2(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT7), .ZN(new_n287));
  XNOR2_X1  g086(.A(G99gat), .B(G106gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G99gat), .A2(G106gat), .ZN(new_n289));
  INV_X1    g088(.A(G85gat), .ZN(new_n290));
  INV_X1    g089(.A(G92gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(KEYINPUT8), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n287), .B2(new_n292), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n285), .A2(new_n295), .B1(KEYINPUT41), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT17), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n298), .A3(new_n284), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n283), .B2(new_n284), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G190gat), .B(G218gat), .Z(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT102), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n296), .A2(KEYINPUT41), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT101), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n307), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n305), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT105), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n218), .A2(new_n219), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n226), .A2(KEYINPUT99), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n293), .A2(KEYINPUT103), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n223), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n295), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n222), .B1(new_n218), .B2(new_n219), .ZN(new_n321));
  INV_X1    g120(.A(new_n295), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(new_n317), .A3(new_n322), .A4(new_n318), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT10), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT104), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n228), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n327), .A3(new_n317), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT104), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n315), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n314), .A3(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G120gat), .B(G148gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G176gat), .B(G204gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n269), .A2(new_n272), .A3(new_n312), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT95), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346));
  INV_X1    g145(.A(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G113gat), .ZN(new_n348));
  INV_X1    g147(.A(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G120gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT1), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n232), .A2(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(G134gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G127gat), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT68), .B1(new_n232), .B2(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n354), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT68), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n356), .B1(new_n359), .B2(new_n351), .ZN(new_n360));
  NOR3_X1   g159(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G148gat), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n361), .A2(new_n363), .B1(new_n365), .B2(KEYINPUT76), .ZN(new_n366));
  INV_X1    g165(.A(G148gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G141gat), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT76), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT2), .B1(new_n365), .B2(new_n368), .ZN(new_n370));
  INV_X1    g169(.A(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n265), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n362), .ZN(new_n373));
  OAI22_X1  g172(.A1(new_n366), .A2(new_n369), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n346), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n265), .A3(new_n371), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n367), .A2(G141gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n377), .A2(new_n362), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT76), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n364), .A2(G148gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n376), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n372), .A2(new_n362), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n380), .A2(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n352), .B2(new_n354), .ZN(new_n387));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n387), .A2(new_n357), .B1(KEYINPUT1), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n389), .A4(new_n356), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT77), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n374), .A2(KEYINPUT3), .B1(new_n389), .B2(new_n356), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n375), .A2(new_n390), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n393), .B1(new_n385), .B2(new_n394), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n378), .A2(new_n379), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n381), .B(new_n404), .C1(new_n363), .C2(new_n361), .ZN(new_n405));
  XNOR2_X1  g204(.A(G141gat), .B(G148gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n362), .B(new_n372), .C1(new_n406), .C2(KEYINPUT2), .ZN(new_n407));
  AND4_X1   g206(.A1(new_n393), .A2(new_n405), .A3(new_n394), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n397), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n402), .A2(new_n409), .A3(new_n399), .A4(new_n400), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n409), .A3(new_n400), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n360), .B(new_n374), .ZN(new_n414));
  INV_X1    g213(.A(new_n400), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n399), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n401), .A2(new_n412), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT0), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  NOR2_X1   g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n414), .A2(new_n415), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI221_X1 g225(.A(new_n426), .B1(new_n425), .B2(new_n424), .C1(new_n400), .C2(new_n398), .ZN(new_n427));
  OR3_X1    g226(.A1(new_n398), .A2(KEYINPUT39), .A3(new_n400), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n428), .A2(new_n429), .A3(new_n421), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n428), .B2(new_n421), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n422), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G211gat), .B(G218gat), .Z(new_n435));
  XOR2_X1   g234(.A(G197gat), .B(G204gat), .Z(new_n436));
  AOI21_X1  g235(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n435), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT72), .B(new_n441), .C1(new_n436), .C2(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT73), .Z(new_n445));
  INV_X1    g244(.A(G183gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT27), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G183gat), .ZN(new_n449));
  INV_X1    g248(.A(G190gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT65), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT28), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT66), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n446), .A2(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(G169gat), .ZN(new_n456));
  INV_X1    g255(.A(G176gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT67), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n456), .A3(new_n457), .A4(KEYINPUT67), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n455), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n451), .B2(KEYINPUT65), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n454), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n450), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G190gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT23), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G169gat), .B2(G176gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(G169gat), .A2(G176gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n473), .A2(new_n475), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT25), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n480), .C1(new_n472), .C2(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n445), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n444), .B1(new_n467), .B2(new_n485), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT74), .B(new_n443), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n445), .ZN(new_n491));
  INV_X1    g290(.A(new_n443), .ZN(new_n492));
  INV_X1    g291(.A(new_n444), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT29), .B1(new_n467), .B2(new_n485), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n486), .A2(new_n493), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n445), .B2(new_n494), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT74), .B1(new_n498), .B2(new_n443), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n501));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(G64gat), .B(G92gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n487), .ZN(new_n507));
  INV_X1    g306(.A(new_n445), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n489), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(new_n492), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(new_n495), .A3(new_n490), .A4(new_n504), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT30), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n496), .B2(new_n499), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n495), .A4(new_n490), .ZN(new_n516));
  INV_X1    g315(.A(new_n504), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n434), .B(new_n519), .C1(new_n433), .C2(new_n432), .ZN(new_n520));
  XNOR2_X1  g319(.A(G78gat), .B(G106gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G22gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G50gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n438), .A2(new_n435), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n441), .B1(new_n436), .B2(new_n437), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n487), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT3), .B1(new_n527), .B2(KEYINPUT80), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(KEYINPUT80), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n374), .ZN(new_n530));
  NAND2_X1  g329(.A1(G228gat), .A2(G233gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n492), .B1(new_n396), .B2(new_n487), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n440), .A2(new_n487), .A3(new_n442), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n385), .B1(new_n535), .B2(new_n394), .ZN(new_n536));
  OAI211_X1 g335(.A(G228gat), .B(G233gat), .C1(new_n532), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n524), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n537), .A3(new_n524), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n522), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  INV_X1    g341(.A(new_n522), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n542), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n413), .A2(new_n416), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n410), .A2(new_n411), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n410), .A2(new_n411), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n421), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(new_n422), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n417), .A2(new_n550), .A3(new_n421), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n511), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n515), .A2(new_n516), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT37), .ZN(new_n557));
  OR3_X1    g356(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT37), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n558), .A2(KEYINPUT38), .A3(new_n517), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT38), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n491), .B(new_n443), .C1(new_n493), .C2(new_n494), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n561), .B(KEYINPUT37), .C1(new_n509), .C2(new_n443), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n517), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n557), .A2(new_n559), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n520), .B(new_n545), .C1(new_n555), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n486), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n467), .A2(new_n485), .A3(KEYINPUT69), .A4(new_n360), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(G227gat), .A3(G233gat), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT32), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G15gat), .B(G43gat), .Z(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G99gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n571), .B(KEYINPUT32), .C1(new_n573), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(new_n570), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n583));
  NAND2_X1  g382(.A1(G227gat), .A2(G233gat), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n566), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n587), .A2(new_n578), .A3(KEYINPUT71), .A4(new_n580), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n588), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n581), .A2(KEYINPUT70), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n597), .A3(new_n580), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n588), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n591), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT79), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(new_n554), .B2(new_n519), .ZN(new_n603));
  INV_X1    g402(.A(new_n545), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n556), .A2(new_n517), .B1(new_n512), .B2(new_n505), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n606));
  INV_X1    g405(.A(new_n421), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n550), .A3(new_n549), .ZN(new_n609));
  INV_X1    g408(.A(new_n553), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n611), .A3(KEYINPUT79), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n604), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n565), .A2(new_n601), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n593), .A2(new_n604), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n554), .A2(new_n519), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n545), .A2(new_n591), .A3(new_n599), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n605), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT79), .B1(new_n605), .B2(new_n611), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n624), .B2(KEYINPUT83), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT83), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n626), .A3(KEYINPUT35), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n615), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT92), .B1(new_n302), .B2(new_n261), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n261), .A2(new_n285), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n285), .A2(KEYINPUT17), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n299), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n258), .A2(new_n260), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .A4(new_n253), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(KEYINPUT94), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n631), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n634), .A2(new_n253), .A3(new_n283), .A4(new_n284), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n630), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G169gat), .B(G197gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n645), .B(new_n651), .C1(new_n637), .C2(new_n638), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n637), .B2(new_n638), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n640), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n651), .B(KEYINPUT85), .ZN(new_n656));
  INV_X1    g455(.A(new_n639), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n645), .B1(new_n637), .B2(new_n638), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n345), .B1(new_n628), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n545), .A2(new_n591), .A3(new_n599), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n603), .B2(new_n612), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT83), .B1(new_n664), .B2(new_n617), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n627), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n614), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(KEYINPUT95), .A3(new_n660), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n344), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n554), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g471(.A(KEYINPUT95), .B1(new_n668), .B2(new_n660), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n345), .B(new_n661), .C1(new_n667), .C2(new_n614), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n519), .B(new_n343), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G8gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT42), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n670), .A2(new_n519), .A3(new_n678), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n683), .B2(new_n676), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(new_n593), .ZN(new_n691));
  AOI21_X1  g490(.A(G15gat), .B1(new_n670), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n601), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT107), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n692), .B1(new_n670), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g495(.A1(new_n670), .A2(new_n604), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n272), .A2(new_n269), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n342), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n312), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n673), .B2(new_n674), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n703), .A2(G29gat), .A3(new_n611), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n668), .B2(new_n311), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n708), .B(new_n312), .C1(new_n667), .C2(new_n614), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  INV_X1    g510(.A(new_n659), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n640), .A2(new_n652), .A3(new_n654), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n639), .B(KEYINPUT94), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT108), .B(new_n659), .C1(new_n715), .C2(new_n652), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n700), .A3(new_n342), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT109), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n554), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G29gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n705), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n723), .A3(new_n724), .ZN(G1328gat));
  OR3_X1    g524(.A1(new_n703), .A2(G36gat), .A3(new_n605), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n519), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G36gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n693), .A3(new_n720), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT47), .B1(new_n733), .B2(KEYINPUT110), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n593), .A2(G43gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n703), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n733), .B1(KEYINPUT110), .B2(KEYINPUT47), .C1(new_n703), .C2(new_n735), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1330gat));
  OAI21_X1  g538(.A(new_n708), .B1(new_n628), .B2(new_n312), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n668), .A2(KEYINPUT44), .A3(new_n311), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n740), .A2(new_n604), .A3(new_n741), .A4(new_n720), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT111), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n710), .A2(new_n744), .A3(new_n604), .A4(new_n720), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n745), .A3(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n545), .A2(G50gat), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n702), .B(new_n747), .C1(new_n673), .C2(new_n674), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT48), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n742), .A2(G50gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n748), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n751), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G50gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n742), .B2(KEYINPUT111), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n749), .B1(new_n759), .B2(new_n745), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT48), .B1(new_n753), .B2(new_n748), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT112), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(G1331gat));
  NOR4_X1   g562(.A1(new_n718), .A2(new_n700), .A3(new_n311), .A4(new_n342), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n668), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n611), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT113), .B(G57gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1332gat));
  XNOR2_X1  g567(.A(new_n605), .B(KEYINPUT114), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n207), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT49), .B(G64gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT115), .Z(G1333gat));
  NOR3_X1   g574(.A1(new_n765), .A2(G71gat), .A3(new_n593), .ZN(new_n776));
  INV_X1    g575(.A(new_n765), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n693), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(G71gat), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n604), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  INV_X1    g582(.A(new_n700), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n718), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n668), .A2(new_n311), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n668), .A2(KEYINPUT51), .A3(new_n311), .A4(new_n785), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT117), .A3(new_n787), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT118), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n342), .A2(G85gat), .A3(new_n611), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n710), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n718), .A2(new_n784), .A3(new_n342), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n611), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n290), .B2(new_n802), .ZN(G1336gat));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n799), .A2(new_n769), .A3(new_n801), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n291), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n769), .A2(G92gat), .A3(new_n342), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n710), .A2(new_n519), .A3(new_n800), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n790), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n807), .B(KEYINPUT119), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n809), .A2(G92gat), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n806), .A2(new_n808), .B1(new_n812), .B2(new_n804), .ZN(G1337gat));
  NOR3_X1   g612(.A1(new_n593), .A2(new_n342), .A3(G99gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n796), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(G99gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n601), .A3(new_n801), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(G1338gat));
  NAND3_X1  g617(.A1(new_n710), .A2(new_n604), .A3(new_n800), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n819), .B2(G106gat), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n342), .A2(G106gat), .A3(new_n545), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n791), .A2(new_n792), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(KEYINPUT120), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(KEYINPUT120), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n819), .A2(G106gat), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n810), .A2(new_n821), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n320), .A2(new_n323), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n326), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(new_n314), .A3(new_n328), .A4(new_n330), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n332), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(new_n315), .C1(new_n324), .C2(new_n331), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n338), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n340), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n835), .A2(new_n338), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n838), .B2(new_n833), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n714), .A2(new_n840), .A3(new_n716), .ZN(new_n841));
  INV_X1    g640(.A(new_n631), .ZN(new_n842));
  INV_X1    g641(.A(new_n629), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n636), .A2(new_n630), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT121), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(KEYINPUT121), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n643), .A2(new_n630), .A3(new_n642), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT122), .Z(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n650), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n655), .A3(new_n341), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n311), .B1(new_n841), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n713), .B1(new_n650), .B2(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n840), .A3(new_n311), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n700), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n343), .A2(new_n717), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n611), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(new_n620), .A3(new_n769), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n718), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n616), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n769), .A2(new_n554), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n661), .A2(new_n349), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  INV_X1    g667(.A(new_n866), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n869), .B2(new_n342), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n341), .A2(new_n347), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT123), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n860), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n869), .B2(new_n700), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n232), .A3(new_n784), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n869), .B2(new_n312), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n312), .A2(new_n519), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n859), .A2(new_n353), .A3(new_n620), .A4(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n545), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n840), .A2(new_n660), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n852), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n312), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n784), .B1(new_n889), .B2(new_n855), .ZN(new_n890));
  INV_X1    g689(.A(new_n858), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n545), .B1(new_n857), .B2(new_n858), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n865), .A2(new_n693), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n884), .B(G141gat), .C1(new_n896), .C2(new_n661), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n859), .A2(KEYINPUT125), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n601), .A2(new_n604), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n859), .B2(KEYINPUT125), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n661), .A2(G141gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n898), .A2(new_n900), .A3(new_n769), .A4(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n897), .B(new_n902), .C1(KEYINPUT126), .C2(new_n884), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(KEYINPUT126), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n894), .A2(KEYINPUT124), .A3(new_n895), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n718), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(G141gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(new_n884), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n341), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n344), .A2(new_n660), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n890), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n604), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n885), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n862), .A2(new_n886), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT59), .B1(new_n917), .B2(new_n367), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n906), .A2(new_n341), .A3(new_n907), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n367), .A2(KEYINPUT59), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n898), .A2(new_n900), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n769), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n367), .A3(new_n341), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n265), .A3(new_n784), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n907), .ZN(new_n927));
  OAI21_X1  g726(.A(G155gat), .B1(new_n927), .B2(new_n700), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n927), .B2(new_n312), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n922), .A2(new_n371), .A3(new_n879), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n554), .A2(new_n605), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n862), .A2(new_n616), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n456), .A3(new_n661), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n554), .B(new_n769), .C1(new_n857), .C2(new_n858), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n620), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n718), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n939), .B2(new_n456), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n934), .B2(new_n342), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n341), .A2(new_n457), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n937), .B2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n934), .B2(new_n700), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n447), .A2(new_n449), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n784), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n937), .A2(KEYINPUT127), .A3(new_n947), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n934), .B2(new_n312), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n450), .A3(new_n311), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  AND3_X1   g758(.A1(new_n936), .A2(new_n604), .A3(new_n601), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n718), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n915), .A2(new_n916), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n601), .A2(new_n933), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n660), .A2(G197gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  OAI21_X1  g766(.A(G204gat), .B1(new_n964), .B2(new_n342), .ZN(new_n968));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n969), .A3(new_n341), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(G1353gat));
  INV_X1    g772(.A(G211gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n960), .A2(new_n974), .A3(new_n784), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT57), .B1(new_n913), .B2(new_n604), .ZN(new_n976));
  INV_X1    g775(.A(new_n916), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n784), .B(new_n963), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  OAI21_X1  g780(.A(G218gat), .B1(new_n964), .B2(new_n312), .ZN(new_n982));
  INV_X1    g781(.A(G218gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n983), .A3(new_n311), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1355gat));
endmodule


