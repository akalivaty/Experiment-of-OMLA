//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n202), .A2(G77), .A3(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n208), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n205), .A2(G50), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n223), .B1(new_n204), .B2(new_n224), .C1(new_n225), .C2(new_n208), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n216), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n217), .A2(new_n218), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n222), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  OAI21_X1  g0051(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n255), .A3(G274), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n258), .B(new_n209), .C1(G41), .C2(G45), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n256), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(new_n228), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n262), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n273), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G58), .A2(G68), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n210), .B1(new_n201), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n210), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n210), .A2(new_n265), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n279), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n210), .A3(G1), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n279), .ZN(new_n290));
  INV_X1    g0090(.A(G50), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n209), .B2(G20), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n290), .A2(new_n292), .B1(new_n291), .B2(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n275), .A2(G169), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n277), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n298), .B(new_n300), .C1(new_n301), .C2(new_n275), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n275), .A2(G190), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n298), .A2(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .A4(new_n303), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n297), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n256), .B1(new_n260), .B2(new_n229), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n312), .B1(new_n230), .B2(new_n267), .C1(new_n270), .C2(new_n224), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(new_n274), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n282), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n318), .B1(G20), .B2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n283), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n279), .B1(new_n228), .B2(new_n289), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n209), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n290), .A2(G77), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n316), .B(new_n326), .C1(G169), .C2(new_n314), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n313), .A2(new_n274), .ZN(new_n329));
  INV_X1    g0129(.A(new_n311), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(G190), .B2(new_n314), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G274), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n274), .A2(new_n336), .A3(new_n252), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n257), .A2(new_n255), .A3(new_n259), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G238), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT70), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G33), .A3(G97), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n263), .A2(G33), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G226), .A4(new_n268), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n346), .ZN(new_n349));
  INV_X1    g0149(.A(G232), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n349), .A2(new_n350), .A3(new_n268), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n274), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n339), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n283), .A2(new_n228), .B1(new_n210), .B2(G68), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n291), .C2(new_n285), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT11), .A3(new_n279), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n288), .A2(G1), .ZN(new_n365));
  NAND2_X1  g0165(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(G20), .A3(new_n204), .A4(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n367), .B(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n204), .B1(new_n209), .B2(G20), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n290), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT11), .B1(new_n363), .B2(new_n279), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n354), .A2(G190), .A3(new_n356), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n358), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n357), .A2(G169), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n354), .A2(G179), .A3(new_n356), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n357), .A2(new_n381), .A3(G169), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n374), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n335), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT69), .B1(new_n310), .B2(new_n334), .ZN(new_n387));
  INV_X1    g0187(.A(new_n290), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n317), .A2(new_n323), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n365), .A2(G20), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n388), .A2(new_n389), .B1(new_n390), .B2(new_n317), .ZN(new_n391));
  INV_X1    g0191(.A(new_n279), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n210), .B1(new_n205), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n285), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n394), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n280), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n318), .A2(G159), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(KEYINPUT74), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n263), .A2(KEYINPUT73), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n406), .A3(G33), .ZN(new_n407));
  AOI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n345), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n204), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n264), .B1(new_n411), .B2(G33), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT7), .B1(new_n412), .B2(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n403), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n392), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n409), .B1(new_n267), .B2(G20), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n409), .A2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(G33), .B1(new_n404), .B2(new_n406), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(new_n266), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n204), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n416), .B1(new_n421), .B2(new_n403), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n391), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(G223), .A2(G1698), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n261), .B2(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n407), .A3(new_n345), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n255), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n337), .B1(new_n338), .B2(G232), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT76), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n256), .B1(new_n260), .B2(new_n350), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n301), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g0236(.A(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n429), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n423), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G169), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n431), .A2(new_n444), .A3(new_n434), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n436), .A2(new_n315), .A3(new_n429), .A4(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n423), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n445), .A2(new_n446), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n414), .A2(KEYINPUT16), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n422), .A3(new_n279), .ZN(new_n451));
  INV_X1    g0251(.A(new_n391), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n449), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n443), .A2(new_n448), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n386), .A2(new_n387), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n255), .A2(G274), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n209), .A2(G45), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n255), .A2(G250), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G238), .A2(G1698), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n229), .B2(G1698), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n407), .A3(new_n345), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n274), .ZN(new_n474));
  AND4_X1   g0274(.A1(KEYINPUT83), .A2(new_n468), .A3(G190), .A4(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n466), .A2(new_n467), .B1(new_n473), .B2(new_n274), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT83), .B1(new_n476), .B2(new_n301), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(G190), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n320), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(new_n390), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n209), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n392), .A2(new_n390), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n225), .ZN(new_n484));
  OR2_X1    g0284(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT82), .B(new_n210), .C1(new_n344), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n341), .A2(new_n343), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G20), .ZN(new_n491));
  NOR3_X1   g0291(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n412), .A2(new_n210), .A3(G68), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n487), .B1(new_n496), .B2(new_n283), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n481), .B(new_n484), .C1(new_n498), .C2(new_n279), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n279), .ZN(new_n500));
  INV_X1    g0300(.A(new_n481), .ZN(new_n501));
  INV_X1    g0301(.A(new_n483), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n480), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(G169), .B1(new_n468), .B2(new_n474), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n315), .B2(new_n476), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n479), .A2(new_n499), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n229), .A2(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n407), .A2(new_n345), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n345), .A2(new_n346), .A3(G250), .A4(G1698), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT4), .A2(G244), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n345), .A2(new_n346), .A3(new_n513), .A4(new_n268), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT79), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n255), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT5), .B(G41), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n274), .B1(new_n460), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G257), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(G274), .A3(new_n255), .A4(new_n460), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n444), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n460), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n274), .A2(new_n336), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n523), .A2(G257), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n510), .B2(new_n509), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n315), .B(new_n531), .C1(new_n533), .C2(new_n255), .ZN(new_n534));
  INV_X1    g0334(.A(new_n418), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n404), .A2(new_n406), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n265), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(new_n346), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT7), .B1(new_n349), .B2(new_n210), .ZN(new_n539));
  OAI21_X1  g0339(.A(G107), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT6), .A2(G97), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(G107), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n230), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G20), .B1(G77), .B2(new_n318), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n392), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  OR3_X1    g0351(.A1(new_n390), .A2(KEYINPUT78), .A3(G97), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT78), .B1(new_n390), .B2(G97), .ZN(new_n553));
  AOI22_X1  g0353(.A1(G97), .A2(new_n502), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n527), .B(new_n534), .C1(new_n551), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n521), .B2(new_n526), .ZN(new_n557));
  OAI211_X1 g0357(.A(G190), .B(new_n531), .C1(new_n533), .C2(new_n255), .ZN(new_n558));
  INV_X1    g0358(.A(new_n550), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n230), .B1(new_n417), .B2(new_n420), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n279), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n554), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n507), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n210), .B1(new_n496), .B2(G33), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n517), .B2(new_n518), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n278), .A2(new_n273), .B1(G20), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(G20), .B1(new_n265), .B2(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n519), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n570), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(KEYINPUT84), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n390), .A2(new_n569), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n502), .B2(new_n569), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n566), .C1(new_n568), .C2(new_n571), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G257), .A2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n216), .B2(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n407), .A3(new_n345), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n349), .A2(G303), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n255), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n528), .A2(G270), .A3(new_n255), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n525), .ZN(new_n588));
  OAI21_X1  g0388(.A(G169), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n565), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n586), .A2(new_n588), .ZN(new_n592));
  INV_X1    g0392(.A(new_n565), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(G169), .A4(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n586), .A2(new_n588), .A3(new_n315), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n591), .B2(new_n595), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n590), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n592), .A2(new_n437), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(G200), .B2(new_n592), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n581), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n523), .A2(G264), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G250), .A2(G1698), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n215), .B2(G1698), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n412), .A2(new_n605), .B1(G33), .B2(G294), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n525), .B(new_n603), .C1(new_n606), .C2(new_n255), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n407), .A3(new_n345), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G33), .A2(G294), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n255), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n525), .A4(new_n603), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(G169), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n528), .A2(G264), .A3(new_n255), .ZN(new_n616));
  INV_X1    g0416(.A(new_n525), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G179), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n289), .A2(new_n230), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT25), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n230), .B2(new_n483), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT22), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n225), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n407), .A2(new_n210), .A3(new_n345), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n210), .A2(G87), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n349), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n472), .A2(G20), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT23), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n210), .B2(G107), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT24), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n624), .B1(new_n636), .B2(new_n279), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n620), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n618), .B2(G200), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n607), .A2(KEYINPUT88), .A3(new_n301), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(G190), .B1(new_n608), .B2(new_n614), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n458), .A2(new_n564), .A3(new_n602), .A4(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n382), .A2(new_n380), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n381), .B1(new_n357), .B2(G169), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n384), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n328), .B2(new_n376), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n443), .A2(new_n456), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n448), .B(new_n455), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n305), .A2(new_n309), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n297), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n556), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT26), .B1(new_n507), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n301), .B1(new_n468), .B2(new_n474), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT83), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n478), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n481), .B1(new_n498), .B2(new_n279), .ZN(new_n663));
  INV_X1    g0463(.A(new_n484), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n476), .A2(KEYINPUT83), .A3(G190), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n504), .A2(new_n506), .ZN(new_n667));
  AND4_X1   g0467(.A1(KEYINPUT26), .A2(new_n666), .A3(new_n667), .A4(new_n658), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n645), .A2(new_n563), .A3(new_n667), .A4(new_n666), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n637), .B1(new_n615), .B2(new_n619), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n599), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n458), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n657), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n365), .A2(new_n210), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n591), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g0485(.A(new_n599), .B(new_n602), .S(new_n685), .Z(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT89), .B1(new_n686), .B2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(KEYINPUT89), .A3(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n684), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n647), .B1(new_n637), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n639), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n599), .A2(new_n691), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n646), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n639), .A2(new_n684), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  NOR2_X1   g0499(.A1(new_n214), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n493), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n221), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NOR2_X1   g0505(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n691), .B1(new_n706), .B2(new_n708), .C1(new_n669), .C2(new_n674), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n684), .B1(new_n670), .B2(new_n675), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n564), .A2(new_n647), .A3(new_n602), .A4(new_n691), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n521), .A2(new_n526), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n618), .ZN(new_n715));
  INV_X1    g0515(.A(new_n476), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n315), .A3(new_n716), .A4(new_n592), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n611), .A2(new_n616), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n714), .A2(new_n595), .A3(new_n476), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n476), .A2(new_n718), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n714), .A4(new_n595), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n717), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n684), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n712), .B1(new_n713), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n711), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n705), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(KEYINPUT91), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n690), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n288), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n209), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n700), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n689), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n687), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT91), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n686), .A2(G330), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n734), .A2(new_n739), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n273), .B1(G20), .B2(new_n444), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n437), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n210), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n496), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n210), .A2(new_n315), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n437), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n437), .A3(G200), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n753), .A2(new_n291), .B1(new_n755), .B2(new_n230), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(G190), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n749), .B(new_n756), .C1(G68), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT93), .B(G159), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT32), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n764), .A2(KEYINPUT32), .B1(G87), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n750), .A2(new_n759), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n267), .B1(new_n769), .B2(new_n228), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n750), .A2(G190), .A3(new_n301), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(G58), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n758), .A2(new_n765), .A3(new_n768), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n349), .B1(new_n769), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n776), .B(new_n778), .C1(G329), .C2(new_n761), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n752), .A2(G326), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n757), .A2(new_n781), .B1(new_n767), .B2(G303), .ZN(new_n782));
  INV_X1    g0582(.A(new_n748), .ZN(new_n783));
  INV_X1    g0583(.A(new_n755), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n783), .A2(G294), .B1(new_n784), .B2(G283), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n746), .B1(new_n774), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n745), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n214), .A2(new_n412), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  INV_X1    g0594(.A(new_n221), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n459), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n459), .C2(new_n250), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n214), .A2(new_n349), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n569), .B2(new_n214), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n792), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n787), .A2(new_n800), .A3(new_n739), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n790), .B(KEYINPUT94), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n686), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n744), .A2(new_n803), .ZN(G396));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n327), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n691), .B1(new_n322), .B2(new_n325), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(new_n333), .B2(new_n332), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n691), .B(new_n811), .C1(new_n669), .C2(new_n674), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n806), .A2(new_n810), .B1(new_n328), .B2(new_n684), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n710), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n738), .B1(new_n815), .B2(new_n729), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n729), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n745), .A2(new_n788), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n739), .B1(new_n228), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n349), .B1(new_n766), .B2(new_n230), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n769), .A2(new_n569), .B1(new_n760), .B2(new_n777), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G294), .B2(new_n772), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n749), .B1(G283), .B2(new_n757), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n752), .A2(G303), .B1(new_n784), .B2(G87), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n821), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n412), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n784), .A2(G68), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n291), .B2(new_n766), .C1(new_n203), .C2(new_n748), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(G132), .C2(new_n761), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n831));
  INV_X1    g0631(.A(new_n769), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n772), .A2(G143), .B1(new_n832), .B2(new_n763), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(new_n757), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n753), .B2(new_n834), .C1(new_n284), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(KEYINPUT97), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT97), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n745), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n819), .B1(new_n841), .B2(new_n843), .C1(new_n814), .C2(new_n789), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n817), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NAND2_X1  g0646(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n220), .A2(new_n569), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n549), .B2(KEYINPUT35), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n795), .A2(G77), .A3(new_n394), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n201), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n209), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n682), .B(KEYINPUT103), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n423), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n457), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n423), .B1(new_n447), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(KEYINPUT104), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n453), .B1(new_n449), .B2(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n441), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(KEYINPUT104), .A3(KEYINPUT37), .A4(new_n441), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n682), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n415), .B1(KEYINPUT16), .B2(new_n414), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n452), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n457), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n864), .A2(new_n875), .A3(new_n441), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n447), .A2(new_n682), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n873), .A2(new_n877), .B1(new_n423), .B2(new_n440), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n384), .A2(new_n684), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT101), .B1(new_n385), .B2(new_n882), .ZN(new_n883));
  AND4_X1   g0683(.A1(KEYINPUT101), .A2(new_n651), .A3(new_n376), .A4(new_n882), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n383), .A2(new_n377), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n883), .A2(new_n884), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n813), .B1(new_n713), .B2(new_n727), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT40), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n874), .B2(new_n879), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n886), .B(new_n887), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n881), .A2(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT106), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n713), .A2(new_n727), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n458), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(G330), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n652), .A2(new_n691), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n870), .A2(new_n900), .A3(new_n880), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT39), .B1(new_n889), .B2(new_n890), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT105), .B1(new_n881), .B2(KEYINPUT39), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n455), .A2(new_n448), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n859), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n885), .A2(new_n882), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n385), .A2(KEYINPUT101), .A3(new_n882), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n651), .A2(new_n376), .A3(new_n882), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n910), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n806), .A2(new_n684), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n812), .B2(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n917), .A2(KEYINPUT102), .B1(new_n889), .B2(new_n890), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n812), .A2(new_n916), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n886), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n909), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n458), .B(new_n709), .C1(new_n710), .C2(new_n708), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n657), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n898), .A2(new_n927), .B1(new_n209), .B2(new_n735), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n898), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n857), .B1(new_n928), .B2(new_n929), .ZN(G367));
  INV_X1    g0730(.A(new_n694), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n684), .B1(new_n551), .B2(new_n555), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n563), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n658), .A2(new_n684), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT108), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n696), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n944), .A3(new_n696), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT43), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n507), .B1(new_n499), .B2(new_n691), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n667), .A2(new_n499), .A3(new_n691), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n639), .B1(new_n939), .B2(new_n940), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n691), .B1(new_n952), .B2(new_n658), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n946), .A2(new_n947), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(new_n953), .A3(new_n945), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n947), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND4_X1   g0758(.A1(new_n931), .A2(new_n954), .A3(new_n941), .A4(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n954), .A2(new_n958), .B1(new_n931), .B2(new_n941), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n700), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(KEYINPUT109), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT45), .B1(new_n941), .B2(new_n698), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  INV_X1    g0766(.A(new_n698), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n939), .C2(new_n940), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n941), .B2(new_n698), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n939), .A2(KEYINPUT44), .A3(new_n967), .A4(new_n940), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n965), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n963), .B1(new_n973), .B2(new_n694), .ZN(new_n974));
  INV_X1    g0774(.A(new_n696), .ZN(new_n975));
  INV_X1    g0775(.A(new_n695), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n693), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n742), .A2(new_n734), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n741), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n731), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n971), .A2(new_n972), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n964), .A2(new_n968), .ZN(new_n984));
  OAI211_X1 g0784(.A(KEYINPUT109), .B(new_n931), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n982), .B(new_n694), .C1(new_n968), .C2(new_n964), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n974), .A2(new_n981), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n962), .B1(new_n987), .B2(new_n731), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n961), .B1(new_n988), .B2(new_n737), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n791), .B1(new_n213), .B2(new_n320), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n794), .B2(new_n243), .ZN(new_n991));
  INV_X1    g0791(.A(G294), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n835), .A2(new_n992), .B1(new_n753), .B2(new_n777), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G97), .B2(new_n784), .ZN(new_n994));
  INV_X1    g0794(.A(G283), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n748), .A2(new_n230), .B1(new_n769), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n772), .A2(G303), .B1(new_n761), .B2(G317), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT46), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n766), .B2(new_n569), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n767), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n827), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n748), .A2(new_n204), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n203), .B2(new_n766), .C1(new_n835), .C2(new_n762), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G150), .A2(new_n772), .B1(new_n202), .B2(new_n832), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n752), .A2(G143), .B1(new_n784), .B2(G77), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n349), .B1(new_n761), .B2(G137), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n999), .A2(new_n1004), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n739), .B(new_n991), .C1(new_n1013), .C2(new_n745), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n950), .B2(new_n802), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n989), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n978), .A2(new_n979), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n730), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n700), .A3(new_n980), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n693), .A2(new_n802), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n771), .A2(new_n291), .B1(new_n769), .B2(new_n204), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G150), .B2(new_n761), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n827), .B1(G97), .B2(new_n784), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n480), .A2(new_n783), .B1(new_n752), .B2(G159), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n757), .A2(new_n317), .B1(new_n767), .B2(G77), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n412), .B1(G326), .B2(new_n761), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n748), .A2(new_n995), .B1(new_n766), .B2(new_n992), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n772), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n753), .B2(new_n775), .C1(new_n777), .C2(new_n835), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1027), .B1(new_n569), .B2(new_n755), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n745), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n702), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n798), .A2(new_n1039), .B1(new_n230), .B2(new_n214), .ZN(new_n1040));
  XOR2_X1   g0840(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(G50), .B2(new_n282), .ZN(new_n1042));
  AOI21_X1  g0842(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n702), .A3(new_n1043), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1041), .A2(G50), .A3(new_n282), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n794), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n240), .A2(new_n459), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n792), .B1(new_n1048), .B2(KEYINPUT112), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT112), .B2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1038), .A2(new_n738), .A3(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1019), .B1(new_n736), .B2(new_n1017), .C1(new_n1020), .C2(new_n1051), .ZN(G393));
  OAI21_X1  g0852(.A(new_n931), .B1(new_n983), .B2(new_n984), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n986), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n736), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n939), .A2(new_n790), .A3(new_n940), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n794), .A2(new_n247), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n792), .B1(G97), .B2(new_n214), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n739), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G317), .A2(new_n752), .B1(new_n772), .B2(G311), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  AOI22_X1  g0863(.A1(G116), .A2(new_n783), .B1(new_n757), .B2(G303), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT114), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT114), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n349), .B1(new_n760), .B2(new_n775), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n230), .A2(new_n755), .B1(new_n766), .B2(new_n995), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G294), .C2(new_n832), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n753), .A2(new_n284), .B1(new_n396), .B2(new_n771), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n317), .A2(new_n832), .B1(new_n761), .B2(G143), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n748), .A2(new_n228), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n204), .A2(new_n766), .B1(new_n755), .B2(new_n225), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n202), .C2(new_n757), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n412), .A3(new_n1073), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n746), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1061), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1055), .B1(new_n1056), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1054), .A2(new_n980), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n987), .A2(new_n1082), .A3(new_n700), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(G390));
  NAND2_X1  g0884(.A1(new_n920), .A2(new_n899), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n905), .A2(new_n906), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n812), .A2(new_n1087), .A3(new_n916), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n812), .B2(new_n916), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n886), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n881), .A2(new_n899), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n886), .A2(new_n728), .A3(new_n814), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1086), .B(new_n1096), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n737), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n818), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n738), .B1(new_n317), .B2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n771), .A2(new_n569), .B1(new_n760), .B2(new_n992), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n267), .B(new_n1103), .C1(G97), .C2(new_n832), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n767), .A2(G87), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n828), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1074), .B1(G283), .B2(new_n752), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n230), .B2(new_n835), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n767), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g0910(.A(G132), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n267), .B1(new_n771), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G125), .B2(new_n761), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G159), .A2(new_n783), .B1(new_n752), .B2(G128), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT120), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n832), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G137), .A2(new_n757), .B1(new_n202), .B2(new_n784), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1106), .A2(new_n1108), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n745), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n906), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n904), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1124), .B2(new_n789), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n458), .A2(new_n728), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n925), .A2(new_n657), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT117), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n925), .A2(new_n1129), .A3(new_n657), .A4(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n886), .B1(new_n728), .B2(new_n814), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1097), .A2(new_n1132), .B1(KEYINPUT118), .B2(new_n813), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n919), .A2(KEYINPUT115), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n812), .A2(new_n1087), .A3(new_n916), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n728), .A2(new_n1136), .A3(new_n814), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n915), .B1(new_n729), .B2(new_n813), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1096), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1133), .A2(new_n1138), .B1(new_n919), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT119), .B1(new_n1131), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n919), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1139), .A2(new_n1096), .B1(new_n1136), .B2(new_n814), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT119), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n1130), .A4(new_n1128), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1098), .A2(new_n1099), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n700), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1100), .B(new_n1125), .C1(new_n1150), .C2(new_n1153), .ZN(G378));
  NAND2_X1  g0954(.A1(new_n294), .A2(new_n871), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n310), .B(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n788), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n738), .B1(new_n202), .B2(new_n1101), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n412), .A2(G41), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n291), .B1(G33), .B2(G41), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n771), .A2(new_n230), .B1(new_n760), .B2(new_n995), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1006), .B1(new_n228), .B2(new_n766), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n480), .C2(new_n832), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n784), .A2(G58), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n753), .B2(new_n569), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G97), .B2(new_n757), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1169), .A3(new_n1161), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n771), .A2(new_n1173), .B1(new_n769), .B2(new_n834), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G132), .B2(new_n757), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1116), .A2(new_n767), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G150), .A2(new_n783), .B1(new_n752), .B2(G125), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n784), .A2(new_n763), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1172), .B(new_n1184), .C1(new_n1171), .C2(new_n1170), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1160), .B1(new_n1185), .B2(new_n745), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1159), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1158), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n893), .B2(G330), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n888), .A2(new_n881), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n891), .A2(new_n892), .ZN(new_n1191));
  AND4_X1   g0991(.A1(G330), .A2(new_n1190), .A3(new_n1191), .A4(new_n1188), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1189), .A2(new_n1192), .B1(new_n907), .B2(new_n923), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1158), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n652), .B(new_n691), .C1(new_n1122), .C2(new_n904), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n893), .A2(G330), .A3(new_n1188), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n889), .A2(new_n890), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n920), .B2(new_n921), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n917), .A2(KEYINPUT102), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1199), .A2(new_n1200), .B1(new_n908), .B2(new_n859), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1193), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1187), .B1(new_n1203), .B2(new_n736), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1131), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1152), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1193), .A2(new_n1202), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(KEYINPUT57), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n700), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1203), .B1(new_n1206), .B2(new_n1152), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT57), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1205), .B1(new_n1210), .B2(new_n1212), .ZN(G375));
  INV_X1    g1013(.A(KEYINPUT122), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1141), .B2(new_n736), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1146), .A2(KEYINPUT122), .A3(new_n737), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n739), .B1(new_n204), .B2(new_n818), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n349), .B1(new_n771), .B2(new_n995), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n783), .A2(new_n480), .B1(new_n784), .B2(G77), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n496), .B2(new_n766), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G303), .C2(new_n761), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n752), .A2(G294), .B1(new_n832), .B2(G107), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n569), .B2(new_n835), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT123), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n753), .A2(new_n1111), .B1(new_n291), .B2(new_n748), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G159), .B2(new_n767), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n769), .A2(new_n284), .B1(new_n760), .B2(new_n1173), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G137), .B2(new_n772), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n412), .A3(new_n1167), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n757), .B2(new_n1116), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1221), .A2(new_n1224), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1217), .B1(new_n746), .B2(new_n1231), .C1(new_n886), .C2(new_n789), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1215), .A2(new_n1216), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n962), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1149), .B2(new_n1236), .ZN(G381));
  OR2_X1    g1037(.A1(G375), .A2(G378), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G387), .A2(new_n1238), .A3(G381), .A4(new_n1239), .ZN(G407));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(G343), .C2(new_n1238), .ZN(G409));
  XNOR2_X1  g1041(.A(G393), .B(G396), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n989), .A2(G390), .A3(new_n1015), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G390), .B1(new_n989), .B2(new_n1015), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1242), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(G393), .B(G396), .Z(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1243), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G378), .B(new_n1205), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1204), .B1(new_n1211), .B2(new_n1235), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1205), .B1(new_n1256), .B2(new_n962), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1100), .A2(new_n1125), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1153), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1262), .A3(KEYINPUT124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1252), .A2(new_n1255), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n683), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1234), .B1(new_n1151), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1131), .A2(new_n1141), .A3(KEYINPUT60), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n700), .A3(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(G384), .A3(new_n1233), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1269), .B2(new_n1233), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(new_n1265), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1272), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(new_n1274), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1275), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1282));
  XOR2_X1   g1082(.A(new_n1272), .B(new_n1282), .Z(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1251), .B1(new_n1281), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1272), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1273), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1283), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1246), .A2(new_n1250), .A3(new_n1285), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1287), .A2(new_n1297), .ZN(G405));
  NAND2_X1  g1098(.A1(G375), .A2(new_n1262), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1279), .A3(new_n1252), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1252), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1272), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1300), .B(new_n1302), .C1(new_n1303), .C2(new_n1251), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1251), .A2(new_n1303), .ZN(new_n1305));
  XOR2_X1   g1105(.A(new_n1304), .B(new_n1305), .Z(G402));
endmodule


