//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT72), .A3(G101), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n463), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n466), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n475), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n487), .B2(G125), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n481), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n478), .B1(new_n489), .B2(G2105), .ZN(G160));
  AND2_X1   g065(.A1(new_n474), .A2(new_n475), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G2105), .A3(new_n473), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n466), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n476), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(G136), .B2(new_n497), .ZN(G162));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n476), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n487), .A2(new_n466), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  AND4_X1   g081(.A1(G2105), .A2(new_n473), .A3(new_n475), .A4(new_n474), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G126), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT73), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n522), .A2(G88), .A3(new_n523), .A4(new_n512), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n522), .A2(G50), .A3(G543), .A4(new_n523), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n522), .A2(new_n523), .A3(new_n512), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n518), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n531), .B1(new_n528), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n532), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n529), .A2(G81), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n518), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT76), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n518), .B1(new_n563), .B2(KEYINPUT76), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n529), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n531), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n531), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OAI221_X1 g149(.A(new_n572), .B1(new_n528), .B2(new_n573), .C1(new_n574), .C2(new_n531), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(G288));
  NAND4_X1  g152(.A1(new_n522), .A2(G86), .A3(new_n523), .A4(new_n512), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n523), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n582), .A2(new_n583), .A3(G651), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n581), .B2(new_n518), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n518), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT79), .ZN(new_n590));
  AOI22_X1  g165(.A1(G47), .A2(new_n532), .B1(new_n529), .B2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n528), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT80), .B(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n532), .A2(G54), .B1(new_n598), .B2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  MUX2_X1   g178(.A(G301), .B(new_n602), .S(new_n603), .Z(G284));
  MUX2_X1   g179(.A(G301), .B(new_n602), .S(new_n603), .Z(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(new_n602), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(new_n555), .B2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  MUX2_X1   g190(.A(KEYINPUT82), .B(new_n613), .S(new_n615), .Z(G323));
  XOR2_X1   g191(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n617));
  XNOR2_X1  g192(.A(G323), .B(new_n617), .ZN(G282));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n492), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(G135), .B2(new_n497), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(KEYINPUT84), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(KEYINPUT84), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(KEYINPUT17), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n651), .B(new_n652), .C1(new_n647), .C2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n648), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n646), .A3(new_n645), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n647), .A3(new_n645), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n667), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n669), .B(new_n672), .C1(new_n664), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  XOR2_X1   g255(.A(new_n575), .B(KEYINPUT86), .Z(new_n681));
  MUX2_X1   g256(.A(G23), .B(new_n681), .S(G16), .Z(new_n682));
  XOR2_X1   g257(.A(KEYINPUT87), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT33), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n682), .B(new_n684), .Z(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G6), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n586), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT32), .B(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G22), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G166), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT88), .B(G1971), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n685), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n686), .A2(G24), .ZN(new_n698));
  INV_X1    g273(.A(G290), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n686), .ZN(new_n700));
  INV_X1    g275(.A(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  INV_X1    g279(.A(G119), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n466), .A2(G107), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n492), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G131), .B2(new_n497), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n696), .A2(new_n697), .A3(new_n702), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT36), .ZN(new_n714));
  NOR2_X1   g289(.A1(G4), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n610), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT89), .B(G1348), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n497), .A2(G141), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT26), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n722), .A2(new_n723), .B1(G105), .B2(new_n464), .ZN(new_n724));
  INV_X1    g299(.A(G129), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n719), .B(new_n724), .C1(new_n725), .C2(new_n492), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G29), .B2(G32), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n686), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n686), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n730), .A2(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n703), .A2(G35), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT95), .Z(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n703), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT29), .Z(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n740), .A2(new_n741), .B1(G1961), .B2(new_n733), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n718), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n623), .A2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n744), .B(new_n745), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n703), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G139), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n476), .B2(new_n757), .C1(new_n758), .C2(new_n466), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n751), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n752), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n686), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n703), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2084), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n762), .A2(new_n767), .A3(new_n773), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n774), .B1(new_n741), .B2(new_n740), .C1(new_n731), .C2(new_n730), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n703), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n497), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n507), .A2(G128), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n466), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT91), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2067), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n686), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n686), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n686), .A2(G19), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n555), .B2(new_n686), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n703), .A2(G27), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G164), .B2(new_n703), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n786), .A2(new_n790), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n743), .A2(new_n775), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n714), .A2(new_n800), .ZN(G150));
  INV_X1    g376(.A(G150), .ZN(G311));
  NOR2_X1   g377(.A1(new_n602), .A2(new_n611), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT38), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n529), .A2(G93), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT96), .B(G55), .Z(new_n807));
  OAI221_X1 g382(.A(new_n805), .B1(new_n518), .B2(new_n806), .C1(new_n531), .C2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(new_n555), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n804), .B(new_n809), .Z(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n811), .A2(new_n812), .A3(G860), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n808), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  OR2_X1    g391(.A1(new_n813), .A2(new_n816), .ZN(G145));
  XNOR2_X1  g392(.A(new_n623), .B(G160), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G162), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n500), .A2(KEYINPUT98), .A3(new_n502), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT98), .B1(new_n500), .B2(new_n502), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n508), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n784), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n726), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n759), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n728), .B2(new_n759), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n824), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n497), .A2(G142), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n507), .A2(G130), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G118), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n832), .A2(KEYINPUT99), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(KEYINPUT99), .B2(new_n832), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(new_n626), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n709), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n828), .B2(KEYINPUT101), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n820), .B1(new_n829), .B2(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(new_n828), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n842), .B(new_n843), .C1(new_n820), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g421(.A1(new_n808), .A2(new_n603), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n681), .B(G303), .ZN(new_n848));
  XNOR2_X1  g423(.A(G290), .B(G305), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT42), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(KEYINPUT42), .C2(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n614), .B(new_n809), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n607), .A2(new_n595), .A3(new_n599), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n600), .A2(G299), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT41), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n859), .B(KEYINPUT102), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n855), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n847), .B1(new_n865), .B2(new_n603), .ZN(G295));
  OAI21_X1  g441(.A(new_n847), .B1(new_n865), .B2(new_n603), .ZN(G331));
  XOR2_X1   g442(.A(new_n850), .B(KEYINPUT103), .Z(new_n868));
  XNOR2_X1  g443(.A(G301), .B(G168), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n809), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n809), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(KEYINPUT106), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n873), .A3(new_n809), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n858), .A3(new_n857), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n860), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  INV_X1    g454(.A(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n861), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n868), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n868), .A2(new_n882), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT43), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n880), .A2(new_n863), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT108), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n875), .A2(new_n861), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n868), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g468(.A1(KEYINPUT43), .A2(new_n889), .A3(new_n893), .A4(new_n843), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT44), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n885), .B2(new_n887), .ZN(new_n897));
  AND4_X1   g472(.A1(new_n896), .A2(new_n889), .A3(new_n893), .A4(new_n843), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n895), .B1(new_n899), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n823), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT45), .B1(new_n902), .B2(KEYINPUT109), .ZN(new_n903));
  INV_X1    g478(.A(new_n506), .ZN(new_n904));
  INV_X1    g479(.A(G126), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n492), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n503), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n500), .A2(KEYINPUT98), .A3(new_n502), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n910), .A2(KEYINPUT109), .A3(G1384), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n497), .A2(G137), .B1(new_n469), .B2(new_n465), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n487), .A2(KEYINPUT69), .A3(G125), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n480), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(G40), .C1(new_n916), .C2(new_n466), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G1996), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n920), .A3(new_n728), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(G1996), .A3(new_n726), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n784), .B(G2067), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n711), .A3(new_n709), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n784), .A2(G2067), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n919), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n918), .B1(new_n726), .B2(new_n923), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT127), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n918), .A2(new_n920), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT46), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n709), .B(new_n711), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n925), .B1(new_n918), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n918), .A2(new_n701), .A3(new_n699), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT48), .ZN(new_n939));
  AOI211_X1 g514(.A(new_n929), .B(new_n935), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT126), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  AND3_X1   g517(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G303), .A2(G8), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(KEYINPUT110), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n945), .A2(new_n950), .A3(G8), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n823), .A2(new_n952), .A3(new_n901), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n509), .A2(new_n901), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n917), .B1(new_n954), .B2(KEYINPUT50), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G2090), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n823), .A2(KEYINPUT45), .A3(new_n901), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n917), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1971), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n917), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n823), .A2(new_n963), .A3(new_n901), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(G1976), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(G288), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n965), .B(new_n967), .C1(new_n966), .C2(new_n681), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n581), .A2(new_n518), .ZN(new_n969));
  OAI21_X1  g544(.A(G1981), .B1(new_n580), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n586), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n586), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT49), .B(new_n970), .C1(new_n973), .C2(new_n974), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n965), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(G8), .B(new_n964), .C1(new_n681), .C2(new_n966), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT52), .ZN(new_n981));
  AND4_X1   g556(.A1(new_n962), .A2(new_n968), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n943), .A2(new_n944), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n917), .B1(new_n902), .B2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(new_n502), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n491), .A2(G138), .A3(new_n466), .A4(new_n473), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(KEYINPUT4), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n952), .B(new_n901), .C1(new_n987), .C2(new_n906), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n503), .B2(new_n508), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(KEYINPUT114), .A3(new_n952), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n984), .A2(new_n741), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n961), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT115), .B(new_n983), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n994), .B2(new_n995), .ZN(new_n1000));
  INV_X1    g575(.A(new_n983), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n982), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n901), .C1(new_n987), .C2(new_n906), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n991), .A2(KEYINPUT116), .A3(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n959), .B1(new_n910), .B2(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n963), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n789), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n953), .A2(new_n955), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n997), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G168), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n1003), .A2(KEYINPUT63), .A3(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n979), .A2(new_n968), .A3(new_n981), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n995), .B1(G2090), .B2(new_n956), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1001), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT63), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n951), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n973), .A2(new_n974), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G288), .A2(G1976), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT112), .Z(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(new_n979), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n965), .A3(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1016), .A2(new_n1020), .A3(new_n1021), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n570), .B2(KEYINPUT117), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(G299), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT50), .B1(new_n910), .B2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n993), .A2(new_n1033), .A3(new_n963), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n766), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n958), .A2(new_n960), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1039));
  INV_X1    g614(.A(G1348), .ZN(new_n1040));
  INV_X1    g615(.A(G2067), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n823), .A2(new_n963), .A3(new_n901), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n956), .A2(new_n1040), .B1(KEYINPUT118), .B2(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n602), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT61), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1956), .B1(new_n984), .B2(new_n993), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n607), .B(new_n1031), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1037), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1051), .B2(new_n1038), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n956), .A2(new_n1040), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n602), .A2(new_n1044), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT60), .B1(new_n1055), .B2(new_n1045), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1049), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1039), .A3(KEYINPUT61), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n958), .A2(new_n960), .A3(new_n920), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n964), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n554), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n610), .A2(new_n1043), .A3(new_n1066), .A4(new_n1044), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1046), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1003), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n982), .A2(new_n998), .A3(KEYINPUT124), .A4(new_n1002), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n958), .A2(new_n960), .A3(new_n797), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n956), .A2(new_n735), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n917), .B1(new_n902), .B2(new_n959), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n1008), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(G301), .A4(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1076), .A2(new_n1083), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT125), .B1(new_n1085), .B2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  OAI21_X1  g662(.A(G2105), .B1(new_n916), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n489), .A2(KEYINPUT123), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n797), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1090), .A2(new_n913), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n912), .A2(new_n958), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1084), .A2(KEYINPUT54), .A3(new_n1086), .A4(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1085), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT122), .B1(new_n1085), .B2(G171), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1080), .A2(G301), .A3(new_n1093), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT54), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1966), .B1(new_n1082), .B2(new_n1008), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1013), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT119), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1011), .A2(new_n1107), .A3(new_n1013), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n997), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT119), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1114));
  OAI21_X1  g689(.A(G8), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1109), .A2(KEYINPUT120), .A3(G8), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1014), .A2(KEYINPUT51), .A3(new_n1110), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1111), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1030), .B1(new_n1103), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1110), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1125), .B2(KEYINPUT51), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1111), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT62), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n1111), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1100), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G290), .B(new_n701), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n937), .B1(new_n919), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n941), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT126), .B(new_n1136), .C1(new_n1122), .C2(new_n1133), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n940), .B1(new_n1138), .B2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g715(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1142));
  NAND2_X1  g716(.A1(new_n1142), .A2(new_n845), .ZN(new_n1143));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n1143), .ZN(G308));
  OR2_X1    g718(.A1(new_n899), .A2(new_n1143), .ZN(G225));
endmodule


