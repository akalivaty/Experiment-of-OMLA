

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n819), .A2(n821), .ZN(n517) );
  INV_X1 U553 ( .A(KEYINPUT103), .ZN(n733) );
  XNOR2_X1 U554 ( .A(n733), .B(KEYINPUT30), .ZN(n734) );
  XNOR2_X1 U555 ( .A(n735), .B(n734), .ZN(n736) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n740) );
  NAND2_X2 U557 ( .A1(n698), .A2(n781), .ZN(n749) );
  NOR2_X1 U558 ( .A1(G651), .A2(n634), .ZN(n648) );
  INV_X1 U559 ( .A(KEYINPUT68), .ZN(n530) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U561 ( .A1(n644), .A2(G85), .ZN(n519) );
  XOR2_X1 U562 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  XNOR2_X1 U563 ( .A(KEYINPUT69), .B(G651), .ZN(n520) );
  NOR2_X1 U564 ( .A1(n634), .A2(n520), .ZN(n645) );
  NAND2_X1 U565 ( .A1(G72), .A2(n645), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n525) );
  NAND2_X1 U567 ( .A1(n648), .A2(G47), .ZN(n523) );
  NOR2_X1 U568 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n521), .Z(n649) );
  NAND2_X1 U570 ( .A1(G60), .A2(n649), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n524) );
  OR2_X1 U572 ( .A1(n525), .A2(n524), .ZN(G290) );
  NAND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U574 ( .A(n526), .B(KEYINPUT67), .ZN(n891) );
  NAND2_X1 U575 ( .A1(G113), .A2(n891), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n527), .Z(n687) );
  NAND2_X1 U578 ( .A1(G137), .A2(n687), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n531), .B(n530), .ZN(n692) );
  XOR2_X1 U581 ( .A(G2104), .B(KEYINPUT64), .Z(n536) );
  NOR2_X1 U582 ( .A1(G2105), .A2(n536), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT65), .B(n532), .Z(n616) );
  NAND2_X1 U584 ( .A1(G101), .A2(n616), .ZN(n534) );
  INV_X1 U585 ( .A(KEYINPUT66), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U587 ( .A(n535), .B(KEYINPUT23), .ZN(n695) );
  AND2_X1 U588 ( .A1(G2105), .A2(n536), .ZN(n892) );
  NAND2_X1 U589 ( .A1(G125), .A2(n892), .ZN(n693) );
  AND2_X1 U590 ( .A1(n695), .A2(n693), .ZN(n537) );
  AND2_X1 U591 ( .A1(n692), .A2(n537), .ZN(G160) );
  XNOR2_X1 U592 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U593 ( .A(KEYINPUT111), .B(G2446), .Z(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT109), .B(G2451), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U596 ( .A(n540), .B(G2430), .Z(n542) );
  XNOR2_X1 U597 ( .A(G1348), .B(G1341), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n542), .B(n541), .ZN(n546) );
  XOR2_X1 U599 ( .A(G2435), .B(KEYINPUT110), .Z(n544) );
  XNOR2_X1 U600 ( .A(G2438), .B(G2454), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U602 ( .A(n546), .B(n545), .Z(n548) );
  XNOR2_X1 U603 ( .A(G2443), .B(G2427), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n548), .B(n547), .ZN(n549) );
  AND2_X1 U605 ( .A1(n549), .A2(G14), .ZN(G401) );
  NAND2_X1 U606 ( .A1(n644), .A2(G90), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G77), .A2(n645), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT9), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G52), .A2(n648), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n649), .A2(G64), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT70), .B(n555), .Z(n556) );
  NOR2_X1 U614 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  XOR2_X1 U616 ( .A(KEYINPUT4), .B(KEYINPUT78), .Z(n559) );
  NAND2_X1 U617 ( .A1(G89), .A2(n644), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT77), .B(n560), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G76), .A2(n645), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U622 ( .A(n563), .B(KEYINPUT5), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n648), .A2(G51), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G63), .A2(n649), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n566), .Z(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U628 ( .A(n569), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G94), .A2(G452), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT71), .ZN(G173) );
  XOR2_X1 U632 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n572) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n572), .B(n571), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n845) );
  NAND2_X1 U636 ( .A1(n845), .A2(G567), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U638 ( .A1(G68), .A2(n645), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT74), .B(n574), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n644), .A2(G81), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT12), .B(n575), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT13), .B(n578), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n649), .A2(G56), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n579), .Z(n582) );
  NAND2_X1 U646 ( .A1(G43), .A2(n648), .ZN(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(n580), .ZN(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n967) );
  INV_X1 U650 ( .A(G860), .ZN(n622) );
  OR2_X1 U651 ( .A1(n967), .A2(n622), .ZN(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(n644), .A2(G92), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G79), .A2(n645), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n648), .A2(G54), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G66), .A2(n649), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n591), .Z(n592) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(n592), .ZN(n714) );
  INV_X1 U662 ( .A(n714), .ZN(n951) );
  NOR2_X1 U663 ( .A1(n951), .A2(G868), .ZN(n594) );
  INV_X1 U664 ( .A(G868), .ZN(n601) );
  NOR2_X1 U665 ( .A1(n601), .A2(G301), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U667 ( .A1(n648), .A2(G53), .ZN(n596) );
  NAND2_X1 U668 ( .A1(G65), .A2(n649), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n644), .A2(G91), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G78), .A2(n645), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n955) );
  XOR2_X1 U674 ( .A(n955), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U675 ( .A1(G299), .A2(G868), .ZN(n603) );
  NOR2_X1 U676 ( .A1(G286), .A2(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U678 ( .A1(G559), .A2(n622), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT79), .B(n604), .Z(n605) );
  NAND2_X1 U680 ( .A1(n714), .A2(n605), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT80), .ZN(n607) );
  XNOR2_X1 U682 ( .A(KEYINPUT16), .B(n607), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n967), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n714), .A2(G868), .ZN(n608) );
  NOR2_X1 U685 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G111), .A2(n891), .ZN(n612) );
  BUF_X1 U688 ( .A(n687), .Z(n895) );
  NAND2_X1 U689 ( .A1(G135), .A2(n895), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n892), .A2(G123), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT18), .B(n613), .Z(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n618) );
  BUF_X1 U694 ( .A(n616), .Z(n896) );
  NAND2_X1 U695 ( .A1(n896), .A2(G99), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n1019) );
  XNOR2_X1 U697 ( .A(G2096), .B(n1019), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n619), .A2(G2100), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT81), .ZN(G156) );
  NAND2_X1 U700 ( .A1(n714), .A2(G559), .ZN(n621) );
  XOR2_X1 U701 ( .A(n967), .B(n621), .Z(n662) );
  NAND2_X1 U702 ( .A1(n622), .A2(n662), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n648), .A2(G55), .ZN(n624) );
  NAND2_X1 U704 ( .A1(G67), .A2(n649), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n644), .A2(G93), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G80), .A2(n645), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n664) );
  XOR2_X1 U710 ( .A(n629), .B(n664), .Z(G145) );
  NAND2_X1 U711 ( .A1(G49), .A2(n648), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U714 ( .A(KEYINPUT82), .B(n632), .ZN(n633) );
  NOR2_X1 U715 ( .A1(n649), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U718 ( .A1(n644), .A2(G86), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G61), .A2(n649), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n645), .A2(G73), .ZN(n639) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n648), .A2(G48), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U726 ( .A1(n644), .A2(G88), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G75), .A2(n645), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n648), .A2(G50), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G62), .A2(n649), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n653), .A2(n652), .ZN(G166) );
  XOR2_X1 U733 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n655) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n664), .B(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(G305), .B(G166), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U739 ( .A(n659), .B(G290), .Z(n660) );
  XNOR2_X1 U740 ( .A(G288), .B(n660), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G299), .B(n661), .ZN(n913) );
  XNOR2_X1 U742 ( .A(n662), .B(n913), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G868), .ZN(n666) );
  OR2_X1 U744 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n670), .A2(G2072), .ZN(n671) );
  XNOR2_X1 U751 ( .A(KEYINPUT86), .B(n671), .ZN(G158) );
  NAND2_X1 U752 ( .A1(G108), .A2(G120), .ZN(n672) );
  NOR2_X1 U753 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G69), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n674), .B(KEYINPUT88), .ZN(n851) );
  NAND2_X1 U756 ( .A1(n851), .A2(G567), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n675), .B(KEYINPUT89), .ZN(n681) );
  NAND2_X1 U758 ( .A1(G132), .A2(G82), .ZN(n676) );
  XNOR2_X1 U759 ( .A(n676), .B(KEYINPUT22), .ZN(n677) );
  XNOR2_X1 U760 ( .A(KEYINPUT87), .B(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n678), .A2(G96), .ZN(n679) );
  OR2_X1 U762 ( .A1(G218), .A2(n679), .ZN(n852) );
  AND2_X1 U763 ( .A1(G2106), .A2(n852), .ZN(n680) );
  NOR2_X1 U764 ( .A1(n681), .A2(n680), .ZN(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n850) );
  NAND2_X1 U768 ( .A1(n850), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G114), .A2(n891), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G126), .A2(n892), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U772 ( .A(KEYINPUT90), .B(n686), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n896), .A2(G102), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n687), .A2(G138), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U776 ( .A1(n691), .A2(n690), .ZN(G164) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  AND2_X1 U778 ( .A1(n692), .A2(G40), .ZN(n694) );
  AND2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U781 ( .A(KEYINPUT91), .B(n697), .Z(n782) );
  INV_X1 U782 ( .A(n782), .ZN(n698) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n781) );
  NAND2_X1 U784 ( .A1(G8), .A2(n749), .ZN(n819) );
  OR2_X1 U785 ( .A1(G1966), .A2(n819), .ZN(n744) );
  INV_X1 U786 ( .A(KEYINPUT27), .ZN(n700) );
  INV_X1 U787 ( .A(n749), .ZN(n726) );
  NAND2_X1 U788 ( .A1(n726), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n749), .A2(G1956), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT99), .ZN(n705) );
  NOR2_X1 U793 ( .A1(n955), .A2(n705), .ZN(n704) );
  XOR2_X1 U794 ( .A(n704), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U795 ( .A1(n955), .A2(n705), .ZN(n721) );
  INV_X1 U796 ( .A(G1996), .ZN(n927) );
  NOR2_X1 U797 ( .A1(n749), .A2(n927), .ZN(n707) );
  XOR2_X1 U798 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n706) );
  XNOR2_X1 U799 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n749), .A2(G1341), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U802 ( .A1(n967), .A2(n710), .ZN(n715) );
  OR2_X1 U803 ( .A1(n714), .A2(n715), .ZN(n719) );
  INV_X1 U804 ( .A(G2067), .ZN(n928) );
  NOR2_X1 U805 ( .A1(n749), .A2(n928), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n711), .B(KEYINPUT101), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n749), .A2(G1348), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n725) );
  XOR2_X1 U814 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n724) );
  XNOR2_X1 U815 ( .A(n725), .B(n724), .ZN(n730) );
  XOR2_X1 U816 ( .A(G1961), .B(KEYINPUT98), .Z(n974) );
  NAND2_X1 U817 ( .A1(n974), .A2(n749), .ZN(n728) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n931) );
  NAND2_X1 U819 ( .A1(n726), .A2(n931), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n737), .A2(G171), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n743) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n749), .ZN(n745) );
  INV_X1 U824 ( .A(G8), .ZN(n731) );
  NOR2_X1 U825 ( .A1(n745), .A2(n731), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n744), .A2(n732), .ZN(n735) );
  NOR2_X1 U827 ( .A1(G168), .A2(n736), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U830 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n748) );
  AND2_X1 U832 ( .A1(n744), .A2(n748), .ZN(n747) );
  NAND2_X1 U833 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n805) );
  AND2_X1 U835 ( .A1(n805), .A2(n819), .ZN(n759) );
  NAND2_X1 U836 ( .A1(n748), .A2(G286), .ZN(n756) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n819), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n752), .A2(G303), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n753), .B(KEYINPUT104), .ZN(n754) );
  OR2_X1 U842 ( .A1(n731), .A2(n754), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n758) );
  INV_X1 U844 ( .A(KEYINPUT32), .ZN(n757) );
  XNOR2_X1 U845 ( .A(n758), .B(n757), .ZN(n807) );
  NAND2_X1 U846 ( .A1(n759), .A2(n807), .ZN(n764) );
  INV_X1 U847 ( .A(n819), .ZN(n762) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U849 ( .A1(G8), .A2(n760), .ZN(n761) );
  OR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U852 ( .A(KEYINPUT106), .B(n765), .Z(n769) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U854 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  NOR2_X1 U855 ( .A1(n819), .A2(n767), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n804) );
  XNOR2_X1 U857 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G140), .A2(n895), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G104), .A2(n896), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G116), .A2(n891), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G128), .A2(n892), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n779), .ZN(n910) );
  XOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .Z(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT93), .B(n780), .ZN(n838) );
  NOR2_X1 U870 ( .A1(n910), .A2(n838), .ZN(n1014) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT92), .ZN(n840) );
  NAND2_X1 U873 ( .A1(n1014), .A2(n840), .ZN(n835) );
  INV_X1 U874 ( .A(n835), .ZN(n802) );
  NAND2_X1 U875 ( .A1(G129), .A2(n892), .ZN(n785) );
  NAND2_X1 U876 ( .A1(G141), .A2(n895), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n896), .A2(G105), .ZN(n786) );
  XOR2_X1 U879 ( .A(KEYINPUT38), .B(n786), .Z(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n891), .A2(G117), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n890) );
  NAND2_X1 U883 ( .A1(G1996), .A2(n890), .ZN(n791) );
  XNOR2_X1 U884 ( .A(n791), .B(KEYINPUT96), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G131), .A2(n895), .ZN(n793) );
  NAND2_X1 U886 ( .A1(G95), .A2(n896), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U888 ( .A(KEYINPUT95), .B(n794), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G107), .A2(n891), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G119), .A2(n892), .ZN(n795) );
  AND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n909) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n909), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n1013) );
  NAND2_X1 U895 ( .A1(n1013), .A2(n840), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n801), .B(KEYINPUT97), .ZN(n831) );
  OR2_X1 U897 ( .A1(n802), .A2(n831), .ZN(n803) );
  OR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n826) );
  NAND2_X1 U899 ( .A1(G1976), .A2(G288), .ZN(n958) );
  AND2_X1 U900 ( .A1(n805), .A2(n958), .ZN(n806) );
  AND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n811) );
  INV_X1 U902 ( .A(n958), .ZN(n809) );
  NOR2_X1 U903 ( .A1(G1976), .A2(G288), .ZN(n815) );
  NOR2_X1 U904 ( .A1(G1971), .A2(G303), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n815), .A2(n808), .ZN(n962) );
  NOR2_X1 U906 ( .A1(n809), .A2(n962), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT105), .ZN(n820) );
  XOR2_X1 U909 ( .A(G1981), .B(G305), .Z(n948) );
  INV_X1 U910 ( .A(n831), .ZN(n813) );
  AND2_X1 U911 ( .A1(n948), .A2(n813), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n835), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n815), .A2(KEYINPUT33), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n819), .A2(n816), .ZN(n817) );
  OR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n821) );
  AND2_X1 U916 ( .A1(n820), .A2(n517), .ZN(n824) );
  INV_X1 U917 ( .A(n821), .ZN(n822) );
  AND2_X1 U918 ( .A1(n822), .A2(KEYINPUT33), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U921 ( .A(G1986), .B(G290), .ZN(n964) );
  NAND2_X1 U922 ( .A1(n964), .A2(n840), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n843) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n890), .ZN(n1010) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n909), .ZN(n1018) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n829) );
  NOR2_X1 U927 ( .A1(n1018), .A2(n829), .ZN(n830) );
  NOR2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(n832), .Z(n833) );
  NOR2_X1 U930 ( .A1(n1010), .A2(n833), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n837), .B(KEYINPUT108), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n910), .A2(n838), .ZN(n1016) );
  NAND2_X1 U935 ( .A1(n839), .A2(n1016), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n844), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n845), .ZN(G217) );
  INV_X1 U940 ( .A(G661), .ZN(n847) );
  NAND2_X1 U941 ( .A1(G2), .A2(G15), .ZN(n846) );
  NOR2_X1 U942 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT112), .B(n848), .Z(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(G188) );
  XNOR2_X1 U946 ( .A(G120), .B(KEYINPUT113), .ZN(G236) );
  INV_X1 U948 ( .A(G132), .ZN(G219) );
  INV_X1 U949 ( .A(G108), .ZN(G238) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G82), .ZN(G220) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(G2678), .B(G2090), .Z(n856) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1961), .B(G1966), .Z(n862) );
  XNOR2_X1 U964 ( .A(G1981), .B(G1971), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(n863), .B(G2474), .Z(n865) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT41), .B(G1956), .Z(n867) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1976), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n892), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n870), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G112), .A2(n891), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n871), .B(KEYINPUT114), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G136), .A2(n895), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G100), .A2(n896), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U981 ( .A1(n877), .A2(n876), .ZN(G162) );
  XNOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U983 ( .A(n1019), .B(KEYINPUT115), .ZN(n878) );
  XNOR2_X1 U984 ( .A(n879), .B(n878), .ZN(n907) );
  NAND2_X1 U985 ( .A1(n892), .A2(G127), .ZN(n880) );
  XOR2_X1 U986 ( .A(KEYINPUT117), .B(n880), .Z(n882) );
  NAND2_X1 U987 ( .A1(n891), .A2(G115), .ZN(n881) );
  NAND2_X1 U988 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U989 ( .A(n883), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U990 ( .A1(G103), .A2(n896), .ZN(n884) );
  NAND2_X1 U991 ( .A1(n885), .A2(n884), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n895), .A2(G139), .ZN(n886) );
  XOR2_X1 U993 ( .A(KEYINPUT116), .B(n886), .Z(n887) );
  NOR2_X1 U994 ( .A1(n888), .A2(n887), .ZN(n1004) );
  XOR2_X1 U995 ( .A(G160), .B(n1004), .Z(n889) );
  XNOR2_X1 U996 ( .A(n890), .B(n889), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U998 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U999 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n895), .ZN(n898) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n896), .ZN(n897) );
  NAND2_X1 U1002 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1003 ( .A(KEYINPUT45), .B(n899), .Z(n900) );
  NOR2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1005 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1006 ( .A(G164), .B(G162), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1008 ( .A(n907), .B(n906), .Z(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1010 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1012 ( .A(n913), .B(G286), .Z(n915) );
  XNOR2_X1 U1013 ( .A(G171), .B(n951), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(n967), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1018 ( .A(KEYINPUT118), .B(n918), .Z(n919) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n919), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n920) );
  XOR2_X1 U1021 ( .A(KEYINPUT119), .B(n920), .Z(n921) );
  NAND2_X1 U1022 ( .A1(G319), .A2(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(G401), .A2(n922), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1027 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1034) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n1028) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n940) );
  XOR2_X1 U1030 ( .A(G2072), .B(G33), .Z(n925) );
  NAND2_X1 U1031 ( .A1(n925), .A2(G28), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G25), .B(G1991), .ZN(n926) );
  XNOR2_X1 U1033 ( .A(n926), .B(KEYINPUT121), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n927), .B(G32), .ZN(n930) );
  XNOR2_X1 U1035 ( .A(n928), .B(G26), .ZN(n929) );
  NAND2_X1 U1036 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1037 ( .A(G27), .B(n931), .Z(n932) );
  NOR2_X1 U1038 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1039 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(KEYINPUT53), .B(n938), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1043 ( .A(G2084), .B(G34), .Z(n941) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(n941), .ZN(n942) );
  NAND2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(n1028), .B(n944), .ZN(n946) );
  INV_X1 U1047 ( .A(G29), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n947), .ZN(n1003) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1053 ( .A(n950), .B(KEYINPUT57), .ZN(n971) );
  XNOR2_X1 U1054 ( .A(G301), .B(G1961), .ZN(n953) );
  XNOR2_X1 U1055 ( .A(G1348), .B(n951), .ZN(n952) );
  NOR2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1057 ( .A(KEYINPUT122), .B(n954), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n955), .B(G1956), .ZN(n956) );
  XNOR2_X1 U1059 ( .A(n956), .B(KEYINPUT123), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1062 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n1001) );
  INV_X1 U1070 ( .A(G16), .ZN(n999) );
  XNOR2_X1 U1071 ( .A(n974), .B(G5), .ZN(n995) );
  XOR2_X1 U1072 ( .A(G1966), .B(G21), .Z(n985) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1074 ( .A(n975), .B(G4), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1076 ( .A(G1341), .B(G19), .ZN(n976) );
  NOR2_X1 U1077 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(G1956), .ZN(n980) );
  XNOR2_X1 U1080 ( .A(G20), .B(n980), .ZN(n981) );
  NOR2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n983), .ZN(n984) );
  NAND2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n991) );
  XOR2_X1 U1085 ( .A(G1986), .B(G24), .Z(n989) );
  XNOR2_X1 U1086 ( .A(G1976), .B(G23), .ZN(n987) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n986) );
  NOR2_X1 U1088 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1089 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1090 ( .A(n991), .B(n990), .Z(n992) );
  NOR2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1092 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1093 ( .A(n996), .B(KEYINPUT126), .ZN(n997) );
  XOR2_X1 U1094 ( .A(KEYINPUT61), .B(n997), .Z(n998) );
  NAND2_X1 U1095 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1096 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1032) );
  XNOR2_X1 U1098 ( .A(G2072), .B(n1004), .ZN(n1007) );
  XNOR2_X1 U1099 ( .A(G164), .B(G2078), .ZN(n1005) );
  XNOR2_X1 U1100 ( .A(n1005), .B(KEYINPUT120), .ZN(n1006) );
  NAND2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1102 ( .A(n1008), .B(KEYINPUT50), .ZN(n1026) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1105 ( .A(n1011), .B(KEYINPUT51), .ZN(n1012) );
  NOR2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1024) );
  INV_X1 U1107 ( .A(n1014), .ZN(n1015) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(G160), .B(G2084), .Z(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(n1034), .B(n1033), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

