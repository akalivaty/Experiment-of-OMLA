

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U550 ( .A1(n716), .A2(n715), .ZN(n760) );
  BUF_X2 U551 ( .A(n864), .Z(n514) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n537), .Z(n864) );
  NOR2_X2 U553 ( .A1(G2105), .A2(n542), .ZN(n865) );
  AND2_X1 U554 ( .A1(n515), .A2(n519), .ZN(n776) );
  NOR2_X1 U555 ( .A1(n517), .A2(n769), .ZN(n718) );
  NOR2_X1 U556 ( .A1(n788), .A2(G1966), .ZN(n517) );
  NAND2_X1 U557 ( .A1(G8), .A2(n760), .ZN(n788) );
  AND2_X1 U558 ( .A1(n688), .A2(G40), .ZN(n715) );
  NOR2_X2 U559 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  NAND2_X1 U560 ( .A1(n784), .A2(n951), .ZN(n515) );
  NAND2_X1 U561 ( .A1(n516), .A2(n774), .ZN(n784) );
  XNOR2_X1 U562 ( .A(n768), .B(KEYINPUT32), .ZN(n516) );
  NOR2_X1 U563 ( .A1(n771), .A2(n517), .ZN(n772) );
  NOR2_X1 U564 ( .A1(n716), .A2(n518), .ZN(n812) );
  INV_X1 U565 ( .A(n715), .ZN(n518) );
  NOR2_X1 U566 ( .A1(n717), .A2(n788), .ZN(n519) );
  NOR2_X1 U567 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U568 ( .A(KEYINPUT23), .ZN(n540) );
  NOR2_X1 U569 ( .A1(G651), .A2(n625), .ZN(n653) );
  XOR2_X1 U570 ( .A(KEYINPUT7), .B(KEYINPUT79), .Z(n536) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n648) );
  NAND2_X1 U572 ( .A1(n648), .A2(G89), .ZN(n520) );
  XNOR2_X1 U573 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n625) );
  XOR2_X1 U575 ( .A(KEYINPUT66), .B(G651), .Z(n526) );
  NOR2_X1 U576 ( .A1(n625), .A2(n526), .ZN(n646) );
  NAND2_X1 U577 ( .A1(G76), .A2(n646), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n524) );
  XOR2_X1 U579 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n523) );
  XNOR2_X1 U580 ( .A(n524), .B(n523), .ZN(n534) );
  XNOR2_X1 U581 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n653), .A2(G51), .ZN(n525) );
  XNOR2_X1 U583 ( .A(n525), .B(KEYINPUT76), .ZN(n529) );
  NOR2_X1 U584 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n527), .Z(n650) );
  NAND2_X1 U586 ( .A1(G63), .A2(n650), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U588 ( .A(n530), .B(KEYINPUT6), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n536), .B(n535), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G69), .ZN(G235) );
  INV_X1 U595 ( .A(G108), .ZN(G238) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  AND2_X1 U598 ( .A1(G137), .A2(n514), .ZN(n539) );
  INV_X1 U599 ( .A(KEYINPUT65), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n539), .B(n538), .ZN(n548) );
  INV_X1 U601 ( .A(G2104), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G101), .A2(n865), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(n546) );
  AND2_X1 U604 ( .A1(G2105), .A2(G2104), .ZN(n868) );
  NAND2_X1 U605 ( .A1(G113), .A2(n868), .ZN(n544) );
  AND2_X1 U606 ( .A1(n542), .A2(G2105), .ZN(n869) );
  NAND2_X1 U607 ( .A1(G125), .A2(n869), .ZN(n543) );
  AND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n688) );
  BUF_X1 U611 ( .A(n688), .Z(G160) );
  NAND2_X1 U612 ( .A1(n514), .A2(G138), .ZN(n550) );
  INV_X1 U613 ( .A(KEYINPUT93), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n865), .A2(G102), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G114), .A2(n868), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G126), .A2(n869), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n557) );
  XOR2_X1 U622 ( .A(n557), .B(KEYINPUT10), .Z(n912) );
  NAND2_X1 U623 ( .A1(n912), .A2(G567), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  XOR2_X1 U625 ( .A(KEYINPUT14), .B(KEYINPUT73), .Z(n560) );
  NAND2_X1 U626 ( .A1(G56), .A2(n650), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G43), .A2(n653), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT74), .B(n561), .Z(n567) );
  NAND2_X1 U630 ( .A1(n648), .A2(G81), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G68), .A2(n646), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U634 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n942) );
  INV_X1 U637 ( .A(G860), .ZN(n599) );
  OR2_X1 U638 ( .A1(n942), .A2(n599), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G90), .A2(n648), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G77), .A2(n646), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U642 ( .A(KEYINPUT9), .B(n572), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n650), .A2(G64), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n653), .A2(G52), .ZN(n573) );
  AND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n653), .A2(G54), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G66), .A2(n650), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G92), .A2(n648), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G79), .A2(n646), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U655 ( .A(KEYINPUT15), .B(n583), .ZN(n600) );
  INV_X1 U656 ( .A(G868), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n600), .A2(n596), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U659 ( .A1(n653), .A2(G53), .ZN(n586) );
  XNOR2_X1 U660 ( .A(n586), .B(KEYINPUT70), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G65), .A2(n650), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U663 ( .A(KEYINPUT71), .B(n589), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G78), .A2(n646), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(KEYINPUT68), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G91), .A2(n648), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U668 ( .A(KEYINPUT69), .B(n593), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G299) );
  NOR2_X1 U670 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n599), .A2(G559), .ZN(n601) );
  INV_X1 U674 ( .A(n600), .ZN(n941) );
  NAND2_X1 U675 ( .A1(n601), .A2(n941), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n942), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n941), .A2(G868), .ZN(n603) );
  NOR2_X1 U679 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G99), .A2(n865), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT82), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G135), .A2(n514), .ZN(n607) );
  XOR2_X1 U684 ( .A(KEYINPUT81), .B(n607), .Z(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G123), .A2(n869), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT80), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G111), .A2(n868), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n929) );
  XNOR2_X1 U692 ( .A(G2096), .B(n929), .ZN(n616) );
  INV_X1 U693 ( .A(G2100), .ZN(n828) );
  NAND2_X1 U694 ( .A1(n616), .A2(n828), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G559), .A2(n941), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(n942), .ZN(n668) );
  NOR2_X1 U697 ( .A1(n668), .A2(G860), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n653), .A2(G55), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G67), .A2(n650), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G93), .A2(n648), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G80), .A2(n646), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n663) );
  XNOR2_X1 U705 ( .A(n624), .B(n663), .ZN(G145) );
  NAND2_X1 U706 ( .A1(G49), .A2(n653), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G87), .A2(n625), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n650), .A2(n628), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n629) );
  XOR2_X1 U711 ( .A(KEYINPUT83), .B(n629), .Z(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G85), .A2(n648), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G47), .A2(n653), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G60), .A2(n650), .ZN(n634) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(n634), .ZN(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G72), .A2(n646), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U721 ( .A1(n648), .A2(G88), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G62), .A2(n650), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n653), .A2(G50), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT86), .B(n641), .Z(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G75), .A2(n646), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G303) );
  NAND2_X1 U729 ( .A1(n646), .A2(G73), .ZN(n647) );
  XNOR2_X1 U730 ( .A(n647), .B(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G86), .A2(n648), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n649), .B(KEYINPUT84), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G48), .A2(n653), .ZN(n654) );
  XNOR2_X1 U736 ( .A(KEYINPUT85), .B(n654), .ZN(n655) );
  NOR2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(G305) );
  NOR2_X1 U739 ( .A1(G868), .A2(n663), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(KEYINPUT89), .ZN(n671) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n661) );
  XNOR2_X1 U742 ( .A(G288), .B(KEYINPUT88), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n663), .B(n662), .ZN(n665) );
  XOR2_X1 U745 ( .A(G290), .B(G303), .Z(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(n666) );
  INV_X1 U747 ( .A(G299), .ZN(n735) );
  XOR2_X1 U748 ( .A(n666), .B(n735), .Z(n667) );
  XNOR2_X1 U749 ( .A(n667), .B(G305), .ZN(n891) );
  XNOR2_X1 U750 ( .A(n891), .B(n668), .ZN(n669) );
  NAND2_X1 U751 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(G295) );
  XOR2_X1 U753 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n673) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U760 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U763 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G96), .A2(n679), .ZN(n820) );
  NAND2_X1 U765 ( .A1(G2106), .A2(n820), .ZN(n684) );
  NOR2_X1 U766 ( .A1(G237), .A2(G238), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G120), .A2(n680), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n681), .A2(G235), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n682), .B(KEYINPUT91), .ZN(n821) );
  NAND2_X1 U770 ( .A1(G567), .A2(n821), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n684), .A2(n683), .ZN(n822) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n685) );
  XNOR2_X1 U773 ( .A(KEYINPUT92), .B(n685), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n822), .A2(n686), .ZN(n819) );
  NAND2_X1 U775 ( .A1(n819), .A2(G36), .ZN(G176) );
  INV_X1 U776 ( .A(G301), .ZN(G171) );
  INV_X1 U777 ( .A(G303), .ZN(G166) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n716) );
  XNOR2_X1 U779 ( .A(KEYINPUT37), .B(G2067), .ZN(n810) );
  NAND2_X1 U780 ( .A1(G140), .A2(n514), .ZN(n690) );
  NAND2_X1 U781 ( .A1(G104), .A2(n865), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n691), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n869), .A2(G128), .ZN(n692) );
  XNOR2_X1 U785 ( .A(n692), .B(KEYINPUT94), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G116), .A2(n868), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U788 ( .A(KEYINPUT35), .B(n695), .Z(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U790 ( .A(KEYINPUT36), .B(n698), .ZN(n888) );
  NOR2_X1 U791 ( .A1(n810), .A2(n888), .ZN(n925) );
  NAND2_X1 U792 ( .A1(n812), .A2(n925), .ZN(n808) );
  NAND2_X1 U793 ( .A1(G131), .A2(n514), .ZN(n700) );
  NAND2_X1 U794 ( .A1(G95), .A2(n865), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G107), .A2(n868), .ZN(n702) );
  NAND2_X1 U797 ( .A1(G119), .A2(n869), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n881) );
  INV_X1 U800 ( .A(G1991), .ZN(n800) );
  NOR2_X1 U801 ( .A1(n881), .A2(n800), .ZN(n713) );
  NAND2_X1 U802 ( .A1(G141), .A2(n514), .ZN(n706) );
  NAND2_X1 U803 ( .A1(G129), .A2(n869), .ZN(n705) );
  NAND2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n865), .A2(G105), .ZN(n707) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n707), .Z(n708) );
  NOR2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n868), .A2(G117), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n885) );
  AND2_X1 U810 ( .A1(n885), .A2(G1996), .ZN(n712) );
  NOR2_X1 U811 ( .A1(n713), .A2(n712), .ZN(n927) );
  INV_X1 U812 ( .A(n927), .ZN(n714) );
  NAND2_X1 U813 ( .A1(n714), .A2(n812), .ZN(n799) );
  NAND2_X1 U814 ( .A1(n808), .A2(n799), .ZN(n795) );
  NAND2_X1 U815 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U816 ( .A(n946), .ZN(n717) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n760), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n718), .B(KEYINPUT100), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n719), .A2(G8), .ZN(n720) );
  XNOR2_X1 U820 ( .A(n720), .B(KEYINPUT30), .ZN(n721) );
  NOR2_X1 U821 ( .A1(n721), .A2(G168), .ZN(n726) );
  XOR2_X1 U822 ( .A(n760), .B(KEYINPUT96), .Z(n736) );
  XNOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .ZN(n996) );
  NAND2_X1 U824 ( .A1(n736), .A2(n996), .ZN(n723) );
  INV_X1 U825 ( .A(G1961), .ZN(n947) );
  NAND2_X1 U826 ( .A1(n947), .A2(n760), .ZN(n722) );
  NAND2_X1 U827 ( .A1(n723), .A2(n722), .ZN(n729) );
  OR2_X1 U828 ( .A1(n729), .A2(G171), .ZN(n724) );
  XNOR2_X1 U829 ( .A(n724), .B(KEYINPUT101), .ZN(n725) );
  XOR2_X1 U830 ( .A(n727), .B(KEYINPUT31), .Z(n728) );
  XNOR2_X1 U831 ( .A(n728), .B(KEYINPUT102), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n729), .A2(G171), .ZN(n757) );
  XNOR2_X1 U833 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n755) );
  NAND2_X1 U834 ( .A1(G2072), .A2(n736), .ZN(n730) );
  XNOR2_X1 U835 ( .A(n730), .B(KEYINPUT27), .ZN(n732) );
  XNOR2_X1 U836 ( .A(G1956), .B(KEYINPUT97), .ZN(n966) );
  NOR2_X1 U837 ( .A1(n736), .A2(n966), .ZN(n731) );
  NOR2_X1 U838 ( .A1(n732), .A2(n731), .ZN(n734) );
  NOR2_X1 U839 ( .A1(n735), .A2(n734), .ZN(n733) );
  XOR2_X1 U840 ( .A(n733), .B(KEYINPUT28), .Z(n753) );
  NAND2_X1 U841 ( .A1(n735), .A2(n734), .ZN(n751) );
  AND2_X1 U842 ( .A1(n760), .A2(G1348), .ZN(n738) );
  AND2_X1 U843 ( .A1(n736), .A2(G2067), .ZN(n737) );
  NOR2_X1 U844 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U845 ( .A1(n941), .A2(n739), .ZN(n749) );
  NAND2_X1 U846 ( .A1(n941), .A2(n739), .ZN(n747) );
  INV_X1 U847 ( .A(G1996), .ZN(n836) );
  NOR2_X1 U848 ( .A1(n760), .A2(n836), .ZN(n741) );
  XOR2_X1 U849 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n740) );
  XNOR2_X1 U850 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U851 ( .A1(n760), .A2(G1341), .ZN(n742) );
  NAND2_X1 U852 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U853 ( .A1(n942), .A2(n744), .ZN(n745) );
  XOR2_X1 U854 ( .A(KEYINPUT64), .B(n745), .Z(n746) );
  NAND2_X1 U855 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U856 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U857 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U858 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U859 ( .A(n755), .B(n754), .ZN(n756) );
  NAND2_X1 U860 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U861 ( .A1(n759), .A2(n758), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n770), .A2(G286), .ZN(n766) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n760), .ZN(n761) );
  XNOR2_X1 U864 ( .A(KEYINPUT103), .B(n761), .ZN(n764) );
  NOR2_X1 U865 ( .A1(G1971), .A2(n788), .ZN(n762) );
  NOR2_X1 U866 ( .A1(G166), .A2(n762), .ZN(n763) );
  NAND2_X1 U867 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U868 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U869 ( .A1(n767), .A2(G8), .ZN(n768) );
  NAND2_X1 U870 ( .A1(G8), .A2(n769), .ZN(n773) );
  INV_X1 U871 ( .A(n770), .ZN(n771) );
  NAND2_X1 U872 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n777) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n775) );
  NOR2_X1 U875 ( .A1(n777), .A2(n775), .ZN(n951) );
  NOR2_X1 U876 ( .A1(n776), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n777), .A2(KEYINPUT33), .ZN(n778) );
  OR2_X1 U878 ( .A1(n788), .A2(n778), .ZN(n779) );
  XOR2_X1 U879 ( .A(G1981), .B(G305), .Z(n956) );
  NAND2_X1 U880 ( .A1(n779), .A2(n956), .ZN(n780) );
  NOR2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n793) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n782) );
  NAND2_X1 U883 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U884 ( .A1(n784), .A2(n783), .ZN(n785) );
  AND2_X1 U885 ( .A1(n785), .A2(n788), .ZN(n791) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XNOR2_X1 U887 ( .A(n786), .B(KEYINPUT24), .ZN(n787) );
  XNOR2_X1 U888 ( .A(n787), .B(KEYINPUT95), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U890 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U893 ( .A(n796), .B(KEYINPUT104), .ZN(n798) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n953) );
  NAND2_X1 U895 ( .A1(n953), .A2(n812), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n815) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n885), .ZN(n914) );
  INV_X1 U898 ( .A(n799), .ZN(n803) );
  AND2_X1 U899 ( .A1(n800), .A2(n881), .ZN(n928) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U901 ( .A1(n928), .A2(n801), .ZN(n802) );
  NOR2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U903 ( .A1(n914), .A2(n804), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n805) );
  XNOR2_X1 U905 ( .A(KEYINPUT105), .B(n805), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n807), .B(n806), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n810), .A2(n888), .ZN(n934) );
  NAND2_X1 U909 ( .A1(n811), .A2(n934), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U912 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n912), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U915 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  NOR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  XOR2_X1 U922 ( .A(KEYINPUT108), .B(n822), .Z(G319) );
  XOR2_X1 U923 ( .A(KEYINPUT42), .B(G2090), .Z(n824) );
  XNOR2_X1 U924 ( .A(G2078), .B(G2072), .ZN(n823) );
  XNOR2_X1 U925 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U926 ( .A(n825), .B(G2096), .Z(n827) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2084), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n832) );
  XOR2_X1 U929 ( .A(KEYINPUT43), .B(G2678), .Z(n830) );
  XOR2_X1 U930 ( .A(KEYINPUT109), .B(n828), .Z(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U932 ( .A(n832), .B(n831), .Z(G227) );
  XOR2_X1 U933 ( .A(KEYINPUT110), .B(G1981), .Z(n834) );
  XOR2_X1 U934 ( .A(G1966), .B(n947), .Z(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n835), .B(KEYINPUT41), .Z(n838) );
  XOR2_X1 U937 ( .A(n836), .B(G1991), .Z(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1956), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U943 ( .A(KEYINPUT111), .B(G2474), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U945 ( .A1(n869), .A2(G124), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U947 ( .A1(G136), .A2(n514), .ZN(n846) );
  NAND2_X1 U948 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U949 ( .A(KEYINPUT112), .B(n848), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G100), .A2(n865), .ZN(n850) );
  NAND2_X1 U951 ( .A1(G112), .A2(n868), .ZN(n849) );
  NAND2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U953 ( .A1(n852), .A2(n851), .ZN(G162) );
  XNOR2_X1 U954 ( .A(G164), .B(G160), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(G162), .ZN(n878) );
  NAND2_X1 U956 ( .A1(G118), .A2(n868), .ZN(n863) );
  NAND2_X1 U957 ( .A1(n869), .A2(G130), .ZN(n854) );
  XNOR2_X1 U958 ( .A(KEYINPUT113), .B(n854), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n865), .A2(G106), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n855), .B(KEYINPUT114), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G142), .A2(n514), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U963 ( .A(KEYINPUT45), .B(n858), .ZN(n859) );
  XNOR2_X1 U964 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  NOR2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n876) );
  NAND2_X1 U967 ( .A1(G139), .A2(n514), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G103), .A2(n865), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G115), .A2(n868), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G127), .A2(n869), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT117), .B(n872), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n873), .ZN(n874) );
  NOR2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n918) );
  XNOR2_X1 U976 ( .A(n876), .B(n918), .ZN(n877) );
  XOR2_X1 U977 ( .A(n878), .B(n877), .Z(n887) );
  XNOR2_X1 U978 ( .A(n929), .B(KEYINPUT118), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n879), .B(KEYINPUT48), .ZN(n880) );
  XOR2_X1 U980 ( .A(n880), .B(KEYINPUT116), .Z(n883) );
  XNOR2_X1 U981 ( .A(n881), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n942), .B(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(G301), .B(n941), .Z(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(G286), .B(n894), .Z(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U992 ( .A(KEYINPUT107), .B(G2427), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2435), .B(G2438), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n904) );
  XOR2_X1 U995 ( .A(G2443), .B(G2451), .Z(n899) );
  XNOR2_X1 U996 ( .A(G2454), .B(G2446), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n900), .B(G2430), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(n905), .A2(G14), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(n911), .A2(G319), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G120), .ZN(G236) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  INV_X1 U1012 ( .A(n912), .ZN(G223) );
  XOR2_X1 U1013 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1015 ( .A(KEYINPUT121), .B(n915), .Z(n916) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n916), .Z(n923) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n917) );
  XNOR2_X1 U1018 ( .A(KEYINPUT122), .B(n917), .ZN(n920) );
  XOR2_X1 U1019 ( .A(G2072), .B(n918), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n921), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n937) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n930), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT120), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n1008) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n1008), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1017) );
  XOR2_X1 U1036 ( .A(KEYINPUT56), .B(G16), .Z(n965) );
  XOR2_X1 U1037 ( .A(n941), .B(G1348), .Z(n944) );
  XNOR2_X1 U1038 ( .A(n942), .B(G1341), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n955) );
  NAND2_X1 U1040 ( .A1(G1971), .A2(G303), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1042 ( .A(n947), .B(G301), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n962) );
  XOR2_X1 U1047 ( .A(G299), .B(G1956), .Z(n960) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(KEYINPUT57), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(KEYINPUT124), .B(n963), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n1014) );
  XOR2_X1 U1055 ( .A(G1961), .B(G5), .Z(n986) );
  XOR2_X1 U1056 ( .A(G1966), .B(G21), .Z(n976) );
  XNOR2_X1 U1057 ( .A(G20), .B(n966), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G6), .B(G1981), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G4), .B(G1348), .Z(n971) );
  XNOR2_X1 U1063 ( .A(KEYINPUT59), .B(n971), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT60), .B(n974), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n984) );
  XOR2_X1 U1067 ( .A(G1986), .B(G24), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT125), .B(n981), .Z(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n987), .B(KEYINPUT126), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n988), .B(KEYINPUT61), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n989), .ZN(n1011) );
  XOR2_X1 U1079 ( .A(G25), .B(G1991), .Z(n990) );
  NAND2_X1 U1080 ( .A1(n990), .A2(G28), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G26), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G2072), .B(G33), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT123), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(n996), .B(G27), .Z(n998) );
  XNOR2_X1 U1087 ( .A(G1996), .B(G32), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(KEYINPUT53), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(G2084), .B(G34), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT54), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G35), .B(G2090), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(G29), .A2(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(G11), .A2(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1018), .ZN(G150) );
  INV_X1 U1104 ( .A(G150), .ZN(G311) );
endmodule

