//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT22), .ZN(new_n204));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT22), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(G141gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT72), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G155gat), .B(G162gat), .Z(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n228));
  OAI21_X1  g027(.A(G141gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n214), .A2(G148gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n221), .A2(new_n223), .A3(new_n226), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n214), .A2(G148gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n220), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(G141gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT70), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n226), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n222), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n213), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(KEYINPUT78), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n213), .B2(new_n243), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n233), .A2(new_n241), .ZN(new_n247));
  OAI211_X1 g046(.A(G228gat), .B(G233gat), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n244), .A2(KEYINPUT78), .ZN(new_n249));
  OR3_X1    g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(G228gat), .A2(G233gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n212), .B2(KEYINPUT77), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(KEYINPUT77), .B2(new_n206), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n247), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n255), .B2(new_n244), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G78gat), .B(G106gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT31), .ZN(new_n259));
  INV_X1    g058(.A(G50gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT79), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n251), .B1(new_n250), .B2(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  INV_X1    g068(.A(G134gat), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G113gat), .ZN(new_n272));
  INV_X1    g071(.A(G113gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G120gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT1), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(KEYINPUT1), .B(G127gat), .C1(new_n272), .C2(new_n274), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281));
  OAI21_X1  g080(.A(G127gat), .B1(new_n281), .B2(KEYINPUT1), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n282), .A3(G134gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n289));
  AOI21_X1  g088(.A(G190gat), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n285), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(KEYINPUT28), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n289), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT66), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n287), .B2(new_n296), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n307), .A2(new_n303), .A3(KEYINPUT26), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT24), .B1(new_n287), .B2(new_n296), .ZN(new_n314));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n306), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n311), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n312), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n315), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n307), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(KEYINPUT25), .A3(new_n313), .A4(new_n320), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n284), .B1(new_n328), .B2(KEYINPUT67), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT64), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT32), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n331), .A2(KEYINPUT34), .A3(new_n333), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT34), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n329), .B(new_n330), .Z(new_n339));
  INV_X1    g138(.A(new_n333), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n336), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  INV_X1    g142(.A(new_n337), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n335), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT33), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n342), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n342), .B2(new_n345), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n269), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n355), .A2(KEYINPUT35), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n357));
  XOR2_X1   g156(.A(G8gat), .B(G36gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G64gat), .ZN(new_n359));
  INV_X1    g158(.A(G92gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G226gat), .ZN(new_n363));
  INV_X1    g162(.A(G233gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n328), .B2(new_n243), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n302), .A2(new_n309), .B1(new_n322), .B2(new_n326), .ZN(new_n367));
  INV_X1    g166(.A(new_n365), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n212), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n367), .B2(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n328), .A2(new_n365), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n213), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT68), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n213), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n357), .B(new_n362), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n373), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n361), .B(KEYINPUT69), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n361), .B1(new_n379), .B2(new_n376), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G85gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT71), .B(G148gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n220), .B1(new_n391), .B2(G141gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n226), .B1(new_n392), .B2(new_n230), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n232), .A2(new_n223), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n241), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n284), .A3(new_n242), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n279), .A2(new_n283), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n395), .B2(new_n284), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT74), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n400), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n397), .A2(new_n399), .A3(new_n404), .A4(new_n402), .ZN(new_n410));
  INV_X1    g209(.A(new_n399), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n247), .A2(new_n401), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n284), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(KEYINPUT5), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT73), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT73), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n410), .A2(new_n417), .A3(KEYINPUT5), .A4(new_n414), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n390), .B(new_n409), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT75), .B1(new_n419), .B2(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(new_n409), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n389), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT75), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n409), .B1(new_n416), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n389), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n422), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(new_n426), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n428), .A2(new_n425), .A3(new_n389), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n385), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n384), .A2(KEYINPUT80), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n378), .B(new_n437), .C1(new_n382), .C2(new_n383), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n428), .A2(new_n389), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT6), .B1(new_n428), .B2(new_n389), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n433), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n355), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT35), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n356), .A2(new_n435), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n379), .A2(KEYINPUT37), .A3(new_n376), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n361), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n374), .B2(new_n377), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n361), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n383), .B1(new_n456), .B2(KEYINPUT38), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n370), .A2(new_n373), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT38), .B1(new_n458), .B2(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n380), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n444), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n412), .A2(new_n411), .A3(new_n413), .ZN(new_n463));
  INV_X1    g262(.A(new_n408), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n407), .B1(new_n402), .B2(new_n404), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n397), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n462), .B(new_n463), .C1(new_n466), .C2(new_n411), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n462), .A3(new_n411), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n389), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  OR3_X1    g269(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n467), .B2(new_n469), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n439), .A2(new_n442), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n269), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n461), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n353), .B2(new_n354), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n336), .A2(new_n341), .A3(new_n337), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n351), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n342), .A2(new_n345), .A3(new_n352), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT36), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n475), .B(new_n483), .C1(new_n435), .C2(new_n474), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n448), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n486), .A2(G1gat), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n489), .B2(G1gat), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g293(.A1(G29gat), .A2(G36gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n495), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G43gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT15), .B1(new_n506), .B2(G50gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n260), .A2(G43gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n513), .A3(new_n496), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT86), .A4(new_n496), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n509), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n506), .A2(G50gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT84), .B(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(new_n506), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT83), .B(KEYINPUT15), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n519), .B(new_n495), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n494), .B(new_n510), .C1(new_n518), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G50gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n530), .A3(new_n506), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n506), .B2(G50gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n509), .B1(new_n532), .B2(new_n523), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(new_n495), .A3(new_n516), .A4(new_n517), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n494), .B1(new_n534), .B2(new_n510), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n493), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n493), .B1(new_n510), .B2(new_n534), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n510), .B1(new_n518), .B2(new_n525), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT17), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n526), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n537), .B1(new_n545), .B2(new_n493), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n546), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(new_n539), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n543), .B(new_n493), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n539), .B(KEYINPUT89), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT13), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT87), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n542), .A2(new_n547), .A3(new_n559), .A4(new_n551), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT11), .B(G169gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n542), .A2(new_n547), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n554), .B2(new_n555), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n551), .A4(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n542), .A3(new_n551), .A4(new_n547), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT91), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n561), .A2(new_n566), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n202), .B1(new_n485), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(KEYINPUT92), .B(new_n573), .C1(new_n448), .C2(new_n484), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AOI211_X1 g381(.A(new_n492), .B(new_n491), .C1(KEYINPUT21), .C2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n287), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT20), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n586), .A2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n582), .A2(KEYINPUT21), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n207), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT8), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n360), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n601), .B2(new_n604), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G99gat), .B(G106gat), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT94), .B1(new_n603), .B2(new_n360), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(KEYINPUT7), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(G85gat), .B2(G92gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n608), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n616), .B(new_n612), .C1(new_n605), .C2(new_n606), .ZN(new_n618));
  INV_X1    g417(.A(new_n608), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n545), .A2(new_n621), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n617), .A2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n543), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n296), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n621), .B1(new_n527), .B2(new_n535), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n628));
  AND4_X1   g427(.A1(new_n296), .A2(new_n627), .A3(new_n628), .A4(new_n625), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n626), .A2(new_n629), .A3(new_n208), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G190gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n296), .A3(new_n625), .ZN(new_n633));
  AOI21_X1  g432(.A(G218gat), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n599), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n208), .B1(new_n626), .B2(new_n629), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n633), .A3(G218gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(KEYINPUT96), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G134gat), .B(G162gat), .Z(new_n639));
  NOR2_X1   g438(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n598), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n618), .B2(new_n619), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n582), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n621), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n617), .A2(new_n620), .A3(KEYINPUT97), .A4(new_n582), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n648), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n647), .B1(new_n652), .B2(new_n654), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  INV_X1    g459(.A(G176gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n659), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n577), .A2(KEYINPUT98), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n575), .B2(new_n576), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(KEYINPUT75), .B(KEYINPUT6), .C1(new_n428), .C2(new_n389), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n431), .A2(new_n429), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n433), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n440), .B(new_n684), .C1(new_n672), .C2(new_n675), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  NAND2_X1  g485(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n440), .B1(new_n672), .B2(new_n675), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT99), .B1(new_n691), .B2(G8gat), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n690), .A2(new_n693), .A3(new_n488), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n688), .A2(new_n689), .B1(new_n692), .B2(new_n694), .ZN(G1325gat));
  NOR2_X1   g494(.A1(new_n353), .A2(new_n354), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n676), .B2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n483), .B(KEYINPUT100), .Z(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n672), .B2(new_n675), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(G15gat), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n676), .A2(new_n269), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  AND3_X1   g503(.A1(new_n596), .A2(KEYINPUT102), .A3(new_n597), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT102), .B1(new_n596), .B2(new_n597), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n573), .A2(new_n670), .ZN(new_n708));
  INV_X1    g507(.A(new_n644), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n712), .B(new_n269), .C1(new_n681), .C2(new_n385), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT103), .B1(new_n435), .B2(new_n474), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n475), .A2(new_n483), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n448), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT105), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n448), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n711), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n485), .A2(new_n644), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(KEYINPUT44), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n707), .B(new_n708), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n681), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(G29gat), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n598), .A2(new_n644), .A3(new_n669), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT101), .Z(new_n733));
  AND2_X1   g532(.A1(new_n577), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n498), .A3(new_n681), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n499), .A3(new_n439), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n727), .B2(new_n440), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1329gat));
  OAI21_X1  g540(.A(G43gat), .B1(new_n727), .B2(new_n483), .ZN(new_n742));
  INV_X1    g541(.A(new_n696), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n707), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n715), .A2(new_n717), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n715), .A2(new_n717), .A3(new_n716), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n722), .B1(new_n751), .B2(new_n448), .ZN(new_n752));
  INV_X1    g551(.A(new_n723), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n710), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n726), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n747), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n698), .A3(new_n708), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(G43gat), .B1(new_n734), .B2(new_n744), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n746), .B1(new_n758), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g558(.A(KEYINPUT107), .B1(new_n727), .B2(new_n474), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n756), .A2(new_n761), .A3(new_n269), .A4(new_n708), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n762), .A3(new_n521), .ZN(new_n763));
  INV_X1    g562(.A(new_n521), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n734), .A2(new_n764), .A3(new_n269), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n521), .B1(new_n727), .B2(new_n474), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n765), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(G1331gat));
  NOR2_X1   g571(.A1(new_n646), .A2(new_n574), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n670), .B(new_n773), .C1(new_n752), .C2(new_n753), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n728), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n669), .B1(new_n721), .B2(new_n723), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n773), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n440), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n785), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT109), .B(new_n787), .C1(new_n780), .C2(new_n783), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n782), .B1(new_n781), .B2(new_n773), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n779), .A3(new_n785), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n777), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n795), .ZN(G1333gat));
  NAND3_X1  g595(.A1(new_n784), .A2(G71gat), .A3(new_n698), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n774), .A2(new_n743), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n797), .B(new_n798), .C1(G71gat), .C2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(G71gat), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n801), .B(new_n699), .C1(new_n780), .C2(new_n783), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(G71gat), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n269), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  INV_X1    g606(.A(new_n598), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n574), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n720), .A2(new_n644), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n644), .A4(new_n809), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n669), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n681), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n670), .B(new_n809), .C1(new_n724), .C2(new_n726), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n603), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(new_n681), .ZN(G1336gat));
  OAI21_X1  g617(.A(G92gat), .B1(new_n816), .B2(new_n440), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n439), .A2(new_n360), .A3(new_n670), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT110), .Z(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT111), .Z(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n812), .B2(new_n813), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n810), .B2(new_n811), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(new_n829), .B2(new_n821), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n819), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n819), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n828), .A2(new_n832), .A3(new_n834), .ZN(G1337gat));
  AOI21_X1  g634(.A(G99gat), .B1(new_n814), .B2(new_n696), .ZN(new_n836));
  INV_X1    g635(.A(G99gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n816), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n838), .B2(new_n698), .ZN(G1338gat));
  OAI21_X1  g638(.A(G106gat), .B1(new_n816), .B2(new_n474), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n474), .A2(G106gat), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n814), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n670), .B(new_n841), .C1(new_n824), .C2(new_n825), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(G1339gat));
  NOR4_X1   g646(.A1(new_n598), .A2(new_n644), .A3(new_n574), .A4(new_n670), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n655), .A2(new_n656), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n647), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n655), .A2(new_n648), .A3(new_n656), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n851), .ZN(new_n852));
  AOI211_X1 g651(.A(KEYINPUT54), .B(new_n648), .C1(new_n655), .C2(new_n656), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n856), .A3(new_n647), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n857), .B2(new_n664), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n852), .B(KEYINPUT55), .C1(new_n854), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n666), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n666), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n853), .B2(new_n665), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n855), .A3(new_n664), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT55), .B1(new_n866), .B2(new_n852), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n546), .A2(new_n539), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n548), .A2(new_n550), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n565), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n570), .B2(new_n572), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n642), .A2(new_n873), .A3(new_n643), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n859), .A2(new_n862), .A3(new_n666), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n862), .B1(new_n859), .B2(new_n666), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n867), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n642), .A2(new_n873), .A3(new_n643), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n873), .A2(new_n670), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n878), .B2(new_n574), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n875), .B(new_n881), .C1(new_n884), .C2(new_n644), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n848), .B1(new_n885), .B2(new_n707), .ZN(new_n886));
  INV_X1    g685(.A(new_n355), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n728), .A2(new_n439), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n574), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n670), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT117), .B(G120gat), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1341gat));
  AOI21_X1  g694(.A(G127gat), .B1(new_n890), .B2(new_n808), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n890), .A2(new_n747), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(G127gat), .ZN(G1342gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n270), .A3(new_n644), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT56), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n270), .B1(new_n890), .B2(new_n644), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n900), .A2(new_n901), .ZN(G1343gat));
  NAND2_X1  g701(.A1(new_n881), .A2(new_n875), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n877), .A2(new_n867), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n574), .A3(new_n863), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n644), .B1(new_n905), .B2(new_n882), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n707), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n848), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n269), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n888), .A2(new_n483), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n573), .A2(new_n860), .A3(new_n867), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n709), .B1(new_n913), .B2(new_n883), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n875), .A3(new_n881), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n848), .B1(new_n915), .B2(new_n598), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n916), .B2(new_n474), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n911), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n574), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT118), .B1(new_n919), .B2(G141gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT58), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n699), .A2(new_n269), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n889), .A3(new_n886), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n573), .A2(G141gat), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n919), .A2(G141gat), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n921), .B(new_n925), .ZN(G1344gat));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n391), .A3(new_n670), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT119), .Z(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n909), .A2(new_n269), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n474), .A2(KEYINPUT57), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n880), .A2(new_n863), .A3(new_n904), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n561), .A2(new_n566), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n570), .A2(new_n572), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n867), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n860), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n935), .A2(new_n936), .B1(new_n670), .B2(new_n873), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(KEYINPUT120), .C1(new_n937), .C2(new_n644), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n598), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT120), .B1(new_n914), .B2(new_n932), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n908), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n930), .A2(KEYINPUT57), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(new_n669), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n912), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n929), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT59), .B(new_n391), .C1(new_n918), .C2(new_n670), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n928), .B1(new_n946), .B2(new_n947), .ZN(G1345gat));
  AOI21_X1  g747(.A(G155gat), .B1(new_n923), .B2(new_n808), .ZN(new_n949));
  INV_X1    g748(.A(new_n918), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(new_n707), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g751(.A(G162gat), .B1(new_n923), .B2(new_n644), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n950), .A2(new_n225), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n644), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n886), .A2(new_n681), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n887), .A2(new_n440), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G169gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n574), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n681), .A2(new_n440), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n743), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n474), .B1(new_n964), .B2(KEYINPUT121), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n965), .B(new_n886), .C1(KEYINPUT121), .C2(new_n964), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n966), .A2(new_n574), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n961), .B1(new_n967), .B2(new_n960), .ZN(G1348gat));
  NAND3_X1  g767(.A1(new_n966), .A2(G176gat), .A3(new_n670), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n661), .B1(new_n958), .B2(new_n669), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(G1349gat));
  AOI21_X1  g770(.A(new_n287), .B1(new_n966), .B2(new_n747), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n958), .B1(new_n288), .B2(new_n289), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n808), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g774(.A(new_n296), .B1(new_n966), .B2(new_n644), .ZN(new_n976));
  XNOR2_X1  g775(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n296), .A3(new_n644), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1351gat));
  OR3_X1    g779(.A1(new_n922), .A2(KEYINPUT123), .A3(new_n440), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT123), .B1(new_n922), .B2(new_n440), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n981), .A2(new_n956), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g782(.A(KEYINPUT124), .B(G197gat), .Z(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n574), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n698), .A2(new_n963), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n942), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n988), .A2(new_n574), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n989), .B2(new_n985), .ZN(G1352gat));
  NAND3_X1  g789(.A1(new_n983), .A2(new_n663), .A3(new_n670), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  NAND2_X1  g791(.A1(new_n944), .A2(new_n987), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G204gat), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1353gat));
  NAND4_X1  g794(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n808), .A4(new_n987), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT57), .B1(new_n886), .B2(new_n474), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n941), .A2(new_n931), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n808), .A4(new_n987), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n996), .A2(new_n1001), .A3(G211gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT63), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n996), .A2(new_n1001), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n983), .A2(new_n207), .A3(new_n808), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1006), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1354gat));
  AOI21_X1  g811(.A(G218gat), .B1(new_n983), .B2(new_n644), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n644), .A2(G218gat), .ZN(new_n1014));
  XOR2_X1   g813(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  AOI21_X1  g814(.A(new_n1013), .B1(new_n988), .B2(new_n1015), .ZN(G1355gat));
endmodule


