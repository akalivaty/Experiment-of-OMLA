//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1380, new_n1381, new_n1382;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT64), .B1(new_n259), .B2(G274), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n209), .B(G274), .C1(G41), .C2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT64), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G1), .B(G13), .C1(new_n265), .C2(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n264), .B1(G226), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n256), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G190), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(G200), .B2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT10), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n218), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n210), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G58), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n278), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n202), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n278), .B1(G1), .B2(new_n210), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n202), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT68), .B1(new_n295), .B2(KEYINPUT9), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n289), .B2(new_n294), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n274), .A2(new_n275), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n271), .A2(G200), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(new_n298), .C1(new_n272), .C2(new_n271), .ZN(new_n301));
  INV_X1    g0101(.A(new_n296), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n271), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n271), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT8), .B(G58), .Z(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n283), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n278), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n291), .A2(new_n251), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n293), .B2(new_n251), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT66), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n319), .B1(new_n206), .B2(new_n248), .C1(new_n252), .C2(new_n223), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n255), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n264), .B1(G244), .B2(new_n269), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G200), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n318), .B(new_n324), .C1(new_n272), .C2(new_n323), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n317), .B1(new_n323), .B2(new_n305), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n327), .A3(new_n322), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT67), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n329), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT67), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n308), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n260), .A2(new_n263), .B1(new_n268), .B2(new_n223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n249), .ZN(new_n339));
  INV_X1    g0139(.A(G232), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G1698), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n337), .B1(new_n342), .B2(new_n248), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT69), .B1(new_n343), .B2(new_n266), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n339), .B(new_n341), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n336), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT69), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n255), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n335), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n352), .B(new_n335), .C1(new_n344), .C2(new_n350), .ZN(new_n355));
  OAI21_X1  g0155(.A(G169), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(new_n353), .ZN(new_n359));
  INV_X1    g0159(.A(new_n335), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n349), .B1(new_n348), .B2(new_n255), .ZN(new_n361));
  AOI211_X1 g0161(.A(KEYINPUT69), .B(new_n266), .C1(new_n347), .C2(new_n336), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n352), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT14), .A3(G169), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT71), .B1(new_n351), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(new_n369), .A3(KEYINPUT13), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n368), .A2(new_n370), .A3(new_n359), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n358), .A2(new_n366), .B1(new_n371), .B2(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n287), .A2(G50), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n210), .B2(G68), .C1(new_n251), .C2(new_n282), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n374), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT12), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n291), .B2(new_n222), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n293), .A2(new_n222), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT11), .B1(new_n374), .B2(new_n277), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n365), .A2(G200), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n368), .A2(new_n370), .A3(new_n359), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n381), .C1(new_n384), .C2(new_n272), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n334), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n284), .A2(new_n222), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n287), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n265), .ZN(new_n397));
  NAND2_X1  g0197(.A1(KEYINPUT3), .A2(G33), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n210), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n345), .A2(new_n346), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(G20), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n399), .A2(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n394), .B(new_n395), .C1(new_n222), .C2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n397), .A3(new_n398), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n400), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n402), .A2(new_n397), .A3(new_n408), .A4(new_n398), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n393), .B1(new_n410), .B2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n404), .B1(new_n411), .B2(new_n395), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n277), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n281), .A2(new_n285), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n291), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n414), .B2(new_n293), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n338), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n248), .B(new_n418), .C1(G223), .C2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n266), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n260), .A2(new_n263), .B1(new_n268), .B2(new_n340), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n272), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G200), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n421), .B2(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AND4_X1   g0228(.A1(KEYINPUT17), .A2(new_n413), .A3(new_n417), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n416), .B1(new_n412), .B2(new_n277), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT17), .B1(new_n430), .B2(new_n428), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n389), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n422), .A2(G179), .A3(new_n424), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n421), .B2(new_n423), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT18), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  AOI22_X1  g0238(.A1(KEYINPUT72), .A2(new_n405), .B1(new_n399), .B2(new_n400), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n222), .B1(new_n439), .B2(new_n409), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT16), .B1(new_n440), .B2(new_n393), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n278), .B1(new_n441), .B2(new_n404), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n438), .B(new_n435), .C1(new_n442), .C2(new_n416), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n413), .A2(new_n417), .A3(new_n428), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n432), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n388), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT25), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n290), .B2(G107), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n290), .A2(new_n452), .A3(G107), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n209), .A2(G33), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n218), .A2(new_n290), .A3(new_n276), .A4(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n453), .A2(new_n455), .B1(new_n457), .B2(G107), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n210), .B2(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n248), .A2(new_n210), .A3(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n248), .A2(new_n469), .A3(new_n210), .A4(G87), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n277), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n473), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n459), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n255), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n258), .A2(G1), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n255), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n482), .A2(KEYINPUT82), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT82), .B1(new_n482), .B2(new_n486), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n484), .A2(new_n266), .A3(G274), .A4(new_n483), .ZN(new_n490));
  AOI21_X1  g0290(.A(G200), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n482), .A2(new_n486), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT83), .A3(new_n272), .A4(new_n490), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n482), .A2(new_n486), .A3(new_n272), .A4(new_n490), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n477), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n290), .A2(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n457), .B2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n287), .A2(G77), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT6), .B1(new_n207), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G20), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n506), .C1(new_n403), .C2(new_n206), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n277), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT74), .B1(new_n507), .B2(new_n277), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n483), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G257), .A3(new_n266), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT76), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n490), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n514), .B2(new_n490), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT75), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n248), .A2(G244), .A3(new_n249), .A4(new_n522), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT75), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n255), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n519), .A2(new_n327), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n514), .A2(new_n490), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n533), .A3(new_n516), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n305), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n510), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n507), .A2(new_n277), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n277), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n534), .A2(G190), .ZN(new_n542));
  AOI21_X1  g0342(.A(G200), .B1(new_n519), .B2(new_n530), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n500), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n498), .A2(new_n536), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n482), .A2(new_n486), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n482), .A2(new_n486), .A3(KEYINPUT82), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(G179), .A3(new_n490), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G274), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n513), .A2(new_n255), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G169), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n476), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n458), .B1(new_n555), .B2(new_n474), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n209), .A2(G45), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G250), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n255), .A2(new_n559), .B1(new_n551), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g0360(.A(G238), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n561));
  OAI211_X1 g0361(.A(G244), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n255), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n327), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n210), .B1(new_n336), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n224), .A2(new_n205), .A3(new_n206), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n210), .B(G68), .C1(new_n345), .C2(new_n346), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n282), .B2(new_n205), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n277), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n311), .A2(new_n291), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n457), .A2(new_n312), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n566), .B(new_n577), .C1(G169), .C2(new_n565), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n565), .A2(KEYINPUT78), .A3(G190), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT78), .B1(new_n565), .B2(G190), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n573), .A2(new_n277), .B1(new_n291), .B2(new_n311), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n457), .A2(G87), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n565), .C2(new_n426), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n564), .A2(new_n255), .ZN(new_n586));
  INV_X1    g0386(.A(new_n560), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n574), .A2(new_n575), .A3(new_n583), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT77), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n581), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n557), .A2(new_n578), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT79), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n248), .A2(new_n597), .A3(G264), .A4(G1698), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n401), .A2(G303), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n248), .A2(G257), .A3(new_n249), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n255), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n513), .A2(new_n266), .ZN(new_n603));
  INV_X1    g0403(.A(G270), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n490), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G283), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n277), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n277), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n290), .A2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n457), .B2(G116), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n305), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n602), .A2(G179), .A3(new_n606), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n618), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT80), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n607), .A2(new_n619), .A3(new_n625), .A4(KEYINPUT21), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT80), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n605), .B1(new_n601), .B2(new_n255), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G190), .ZN(new_n629));
  INV_X1    g0429(.A(new_n623), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n426), .C2(new_n628), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n624), .A2(new_n626), .A3(new_n627), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n594), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n451), .A2(new_n545), .A3(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n566), .A2(new_n577), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n565), .A2(G169), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n565), .A2(G190), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n635), .A2(new_n636), .B1(new_n584), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT84), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n578), .B(KEYINPUT84), .C1(new_n584), .C2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n498), .A3(new_n536), .A4(new_n544), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n554), .A2(new_n556), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n578), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n510), .A2(new_n531), .A3(new_n535), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT26), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n593), .A2(new_n578), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n536), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n451), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n307), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n413), .A2(new_n417), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n438), .B1(new_n658), .B2(new_n435), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n430), .A2(new_n436), .A3(KEYINPUT18), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n437), .A2(new_n443), .A3(KEYINPUT85), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n329), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n382), .B1(new_n385), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n432), .A2(new_n449), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n656), .B1(new_n667), .B2(new_n304), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n655), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n556), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n498), .A2(new_n557), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n675), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n644), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n677), .A2(new_n679), .B1(new_n645), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n630), .A2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n644), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n632), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT86), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n686), .A3(G330), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n498), .A2(new_n557), .A3(new_n676), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n557), .B2(new_n678), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT87), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n624), .A2(new_n627), .ZN(new_n693));
  INV_X1    g0493(.A(new_n681), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n626), .A3(new_n631), .A4(new_n694), .ZN(new_n695));
  AOI211_X1 g0495(.A(KEYINPUT86), .B(new_n692), .C1(new_n695), .C2(new_n682), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n686), .B1(new_n683), .B2(G330), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT87), .B(new_n690), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n680), .B1(new_n691), .B2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n213), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n569), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n216), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n651), .B1(new_n642), .B2(new_n648), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n650), .A2(new_n536), .A3(KEYINPUT26), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n678), .B1(new_n710), .B2(new_n647), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n678), .C1(new_n647), .C2(new_n653), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n498), .A2(new_n536), .A3(new_n544), .ZN(new_n716));
  NOR4_X1   g0516(.A1(new_n716), .A2(new_n594), .A3(new_n632), .A4(new_n675), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n530), .A2(new_n533), .A3(new_n516), .A4(new_n565), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n602), .A2(new_n606), .A3(G179), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT88), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(KEYINPUT30), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n721), .A2(new_n489), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n724), .B1(new_n721), .B2(new_n489), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT89), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n565), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n534), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n548), .A2(new_n490), .A3(new_n549), .ZN(new_n732));
  AOI21_X1  g0532(.A(G179), .B1(new_n602), .B2(new_n606), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(KEYINPUT90), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n733), .A2(new_n534), .A3(new_n729), .A4(new_n730), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n487), .A2(new_n488), .A3(new_n552), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n727), .A2(new_n739), .A3(KEYINPUT91), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n675), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT91), .B1(new_n727), .B2(new_n739), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n717), .A2(new_n718), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n736), .A2(new_n737), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n718), .B(new_n678), .C1(new_n727), .C2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n692), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n715), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n707), .B1(new_n749), .B2(G1), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT92), .ZN(G364));
  AND2_X1   g0551(.A1(new_n210), .A2(G13), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n209), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n702), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n701), .A2(new_n401), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G355), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G116), .B2(new_n213), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n701), .A2(new_n248), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n258), .B2(new_n217), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n243), .A2(new_n258), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n218), .B1(G20), .B2(new_n305), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n210), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT94), .Z(new_n769));
  OAI21_X1  g0569(.A(new_n755), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n272), .A2(new_n426), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n210), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n772), .A2(new_n272), .A3(G200), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n248), .B1(new_n773), .B2(new_n224), .C1(new_n206), .C2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n272), .A3(new_n426), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n272), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n327), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n205), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT32), .ZN(new_n784));
  INV_X1    g0584(.A(new_n776), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(G159), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n775), .A2(new_n778), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(G20), .A2(G179), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT95), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n789), .A2(KEYINPUT97), .A3(new_n771), .ZN(new_n790));
  AOI21_X1  g0590(.A(KEYINPUT97), .B1(new_n789), .B2(new_n771), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n272), .A3(G200), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n787), .B1(new_n202), .B2(new_n792), .C1(new_n222), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n789), .A2(new_n272), .A3(new_n426), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n789), .A2(new_n779), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n795), .A2(new_n251), .B1(new_n796), .B2(new_n284), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  INV_X1    g0598(.A(new_n774), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G283), .B1(new_n785), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(new_n773), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n248), .B1(new_n801), .B2(G303), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G294), .B2(new_n781), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n795), .C1(new_n792), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n793), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  INV_X1    g0609(.A(new_n796), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n808), .A2(new_n809), .B1(new_n810), .B2(G322), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT98), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n794), .A2(new_n798), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n770), .B1(new_n813), .B2(new_n764), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n767), .B(KEYINPUT99), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n683), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT100), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n695), .A2(new_n692), .A3(new_n682), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n755), .B1(new_n820), .B2(KEYINPUT93), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(KEYINPUT93), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n822), .B2(new_n688), .ZN(G396));
  NAND2_X1  g0623(.A1(new_n329), .A2(KEYINPUT102), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT102), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n326), .A2(new_n825), .A3(new_n328), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n325), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n678), .B(new_n828), .C1(new_n647), .C2(new_n653), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n654), .A2(new_n678), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n317), .A2(new_n678), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n827), .A2(new_n831), .B1(new_n329), .B2(new_n678), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n748), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n755), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n764), .A2(new_n766), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n755), .B1(G77), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G311), .A2(new_n785), .B1(new_n801), .B2(G107), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n401), .C1(new_n224), .C2(new_n774), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n783), .B(new_n841), .C1(G294), .C2(new_n810), .ZN(new_n842));
  INV_X1    g0642(.A(new_n795), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G116), .A2(new_n843), .B1(new_n808), .B2(G283), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n842), .B(new_n844), .C1(new_n845), .C2(new_n792), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT101), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n808), .A2(G150), .B1(new_n810), .B2(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n777), .B2(new_n795), .C1(new_n849), .C2(new_n792), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(KEYINPUT34), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n248), .B1(new_n773), .B2(new_n202), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n774), .A2(new_n222), .B1(new_n776), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G58), .C2(new_n781), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n847), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n839), .B1(new_n859), .B2(new_n764), .ZN(new_n860));
  INV_X1    g0660(.A(new_n766), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n832), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n836), .A2(new_n862), .ZN(G384));
  OR2_X1    g0663(.A1(new_n503), .A2(new_n505), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(G116), .A3(new_n219), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT36), .Z(new_n868));
  OAI211_X1 g0668(.A(new_n217), .B(G77), .C1(new_n284), .C2(new_n222), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n202), .A2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n209), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n430), .A2(new_n673), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n437), .A2(new_n443), .A3(KEYINPUT85), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT85), .B1(new_n437), .B2(new_n443), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n429), .B2(new_n431), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n447), .A2(KEYINPUT105), .A3(new_n448), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n873), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n673), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n442), .B2(new_n416), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n658), .A2(new_n435), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n445), .A4(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n445), .A3(new_n884), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n873), .B2(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n881), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  OR2_X1    g0695(.A1(KEYINPUT103), .A2(KEYINPUT16), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n411), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n277), .B1(new_n411), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n417), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n883), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n435), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n445), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n887), .A2(new_n882), .A3(new_n445), .A4(new_n884), .ZN(new_n904));
  INV_X1    g0704(.A(new_n900), .ZN(new_n905));
  AOI221_X4 g0705(.A(new_n895), .B1(new_n903), .B2(new_n904), .C1(new_n450), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n832), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n381), .A2(new_n678), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n385), .B(new_n910), .C1(new_n372), .C2(new_n381), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n358), .A2(new_n366), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n327), .B2(new_n384), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n909), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n740), .A2(new_n675), .ZN(new_n916));
  INV_X1    g0716(.A(new_n742), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n633), .A2(new_n545), .A3(new_n678), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(KEYINPUT31), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n741), .A2(new_n718), .A3(new_n742), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT40), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n911), .A2(new_n914), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n832), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n917), .A2(KEYINPUT31), .A3(new_n675), .A4(new_n740), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n743), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n450), .A2(new_n905), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n903), .A2(new_n904), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n895), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n926), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n743), .A2(new_n925), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n451), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n692), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n935), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n894), .B2(new_n906), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n382), .A2(new_n678), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n931), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n911), .A2(new_n914), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n824), .A2(new_n826), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n678), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n829), .B2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n932), .A2(new_n949), .B1(new_n876), .B2(new_n673), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n715), .A2(new_n451), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n668), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n939), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n209), .B2(new_n752), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n939), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n872), .B1(new_n956), .B2(new_n957), .ZN(G367));
  OR2_X1    g0758(.A1(new_n590), .A2(new_n678), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n578), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT106), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n642), .A2(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n963), .A2(new_n964), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n815), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n769), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n213), .B2(new_n311), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n760), .A2(new_n239), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n755), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n792), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G143), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n810), .A2(G150), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n782), .A2(new_n222), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n849), .A2(new_n776), .B1(new_n773), .B2(new_n284), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n774), .A2(new_n251), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n978), .A2(new_n401), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G50), .A2(new_n843), .B1(new_n808), .B2(G159), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n976), .A2(new_n977), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n773), .A2(new_n610), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT46), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G107), .B2(new_n781), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT109), .B(G317), .Z(new_n987));
  OAI221_X1 g0787(.A(new_n401), .B1(new_n774), .B2(new_n205), .C1(new_n776), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G303), .B2(new_n810), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G283), .A2(new_n843), .B1(new_n808), .B2(G294), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n792), .A2(new_n805), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n974), .B1(new_n994), .B2(new_n764), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n970), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n749), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n690), .B1(new_n696), .B2(new_n697), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT87), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n648), .A2(new_n675), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n510), .A2(new_n675), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n544), .A2(new_n536), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT45), .B1(new_n680), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n645), .A2(new_n678), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n644), .A2(new_n678), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n689), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1004), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(KEYINPUT44), .A3(new_n1009), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1005), .A2(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1000), .A2(new_n1014), .A3(new_n698), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1000), .B2(new_n698), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n677), .A2(new_n679), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n690), .B2(new_n679), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n688), .B(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n997), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n702), .B(KEYINPUT41), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n753), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n691), .A2(new_n699), .A3(new_n1009), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n967), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT43), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n965), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT42), .B1(new_n1018), .B2(new_n1009), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n536), .B1(new_n1003), .B2(new_n557), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n678), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n689), .A2(new_n1007), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT42), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n1004), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1025), .A2(new_n1028), .A3(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1037), .A2(new_n968), .A3(new_n1027), .A4(new_n1034), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1024), .B(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT108), .B1(new_n1023), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1013), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1008), .A2(KEYINPUT44), .A3(new_n1009), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1010), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1042), .A2(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n691), .B2(new_n699), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1000), .A2(new_n1014), .A3(new_n698), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1047), .A2(new_n749), .A3(new_n1048), .A4(new_n1020), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1022), .B1(new_n1049), .B2(new_n749), .ZN(new_n1050));
  OAI211_X1 g0850(.A(KEYINPUT108), .B(new_n1040), .C1(new_n1050), .C2(new_n754), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n996), .B1(new_n1041), .B2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n1020), .A2(new_n754), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n401), .B1(new_n776), .B2(new_n806), .C1(new_n610), .C2(new_n774), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n808), .A2(G311), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n845), .B2(new_n795), .C1(new_n796), .C2(new_n987), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G322), .B2(new_n975), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n781), .A2(G283), .B1(new_n801), .B2(G294), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1055), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n414), .A2(new_n793), .B1(new_n795), .B2(new_n222), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n782), .A2(new_n311), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n248), .B1(new_n774), .B2(new_n205), .ZN(new_n1068));
  INV_X1    g0868(.A(G150), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1069), .A2(new_n776), .B1(new_n773), .B2(new_n251), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n202), .B2(new_n796), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1066), .B(new_n1072), .C1(G159), .C2(new_n975), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n764), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n755), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n704), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n756), .A2(new_n1076), .B1(new_n206), .B2(new_n701), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n236), .A2(new_n258), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n309), .A2(new_n202), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n704), .B(new_n258), .C1(new_n222), .C2(new_n251), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n759), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1077), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1075), .B1(new_n1083), .B2(new_n971), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1074), .B(new_n1084), .C1(new_n690), .C2(new_n815), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1054), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n749), .A2(new_n1020), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(new_n703), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n749), .A2(new_n1020), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(G393));
  OR2_X1    g0890(.A1(new_n1017), .A2(new_n1087), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n703), .B1(new_n1017), .B2(new_n1087), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n971), .B1(new_n205), .B2(new_n213), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n760), .A2(new_n246), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n755), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n975), .A2(G317), .B1(G311), .B2(new_n810), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G322), .A2(new_n785), .B1(new_n801), .B2(G283), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n248), .B1(new_n799), .B2(G107), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n610), .C2(new_n782), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G303), .B2(new_n808), .ZN(new_n1102));
  INV_X1    g0902(.A(G294), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n795), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n792), .A2(new_n1069), .B1(new_n777), .B2(new_n796), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n808), .A2(G50), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n782), .A2(new_n251), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n401), .B1(new_n799), .B2(G87), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G143), .A2(new_n785), .B1(new_n801), .B2(G68), .ZN(new_n1113));
  AND4_X1   g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1108), .B(new_n1114), .C1(new_n279), .C2(new_n795), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1098), .A2(new_n1104), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1096), .B1(new_n1116), .B2(new_n764), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n767), .B2(new_n1004), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1017), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1093), .B(new_n1118), .C1(new_n1119), .C2(new_n753), .ZN(G390));
  AND3_X1   g0920(.A1(new_n936), .A2(G330), .A3(new_n915), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n829), .A2(new_n948), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n923), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n941), .A2(new_n944), .B1(new_n1123), .B2(new_n942), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n678), .B(new_n828), .C1(new_n710), .C2(new_n647), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n946), .B1(new_n1125), .B2(new_n948), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n907), .A2(new_n1126), .A3(new_n943), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1121), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n878), .A2(new_n879), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n884), .B1(new_n1129), .B2(new_n663), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n895), .B1(new_n1130), .B2(new_n892), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT39), .B1(new_n1131), .B2(new_n931), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT38), .B1(new_n927), .B2(new_n928), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n906), .A2(new_n1133), .A3(new_n940), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1132), .A2(new_n1134), .B1(new_n943), .B2(new_n949), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n915), .B(G330), .C1(new_n919), .C2(new_n746), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n931), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n948), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n942), .B(new_n1137), .C1(new_n1139), .C2(new_n946), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n692), .B1(new_n743), .B2(new_n925), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n451), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n952), .A2(new_n1144), .A3(new_n668), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n832), .C1(new_n919), .C2(new_n746), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n946), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n915), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1147), .A2(new_n1148), .B1(new_n829), .B2(new_n948), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n923), .B1(new_n1143), .B2(new_n832), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1145), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1142), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n923), .B1(new_n748), .B2(new_n832), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1122), .B1(new_n1155), .B2(new_n1121), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n692), .B(new_n908), .C1(new_n743), .C2(new_n925), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1139), .B(new_n1136), .C1(new_n1157), .C2(new_n923), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(new_n1128), .A3(new_n1141), .A4(new_n1145), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n702), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1128), .A2(new_n1141), .A3(new_n754), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n766), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n796), .A2(new_n854), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n801), .A2(G150), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G159), .C2(new_n781), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n248), .B1(new_n776), .B2(new_n1168), .C1(new_n202), .C2(new_n774), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(KEYINPUT111), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G137), .B2(new_n808), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT54), .B(G143), .Z(new_n1172));
  AOI22_X1  g0972(.A1(new_n1169), .A2(KEYINPUT111), .B1(new_n843), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n975), .A2(G128), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1167), .A2(new_n1171), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n975), .A2(G283), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n810), .A2(G116), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n401), .B1(new_n773), .B2(new_n224), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n774), .A2(new_n222), .B1(new_n776), .B2(new_n1103), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1110), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G97), .A2(new_n843), .B1(new_n808), .B2(G107), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n765), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1075), .B(new_n1183), .C1(new_n414), .C2(new_n837), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1163), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1162), .A2(KEYINPUT112), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT112), .B1(new_n1162), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1161), .B1(new_n1186), .B2(new_n1187), .ZN(G378));
  AOI21_X1  g0988(.A(new_n933), .B1(new_n926), .B2(new_n1137), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n933), .B1(new_n906), .B2(new_n1133), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(new_n921), .ZN(new_n1191));
  OAI21_X1  g0991(.A(G330), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n295), .A2(new_n673), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n308), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n308), .A2(new_n1193), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OR3_X1    g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n945), .A2(new_n950), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n945), .B2(new_n950), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1192), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n951), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n692), .B1(new_n922), .B2(new_n934), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n945), .A2(new_n950), .A3(new_n1200), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n766), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n755), .B1(G50), .B2(new_n838), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G50), .B1(new_n398), .B2(new_n257), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G41), .B(new_n248), .C1(new_n801), .C2(G77), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n799), .A2(G58), .B1(new_n785), .B2(G283), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n206), .C2(new_n796), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G97), .B2(new_n808), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n978), .B1(new_n975), .B2(G116), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT113), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1216), .B1(new_n311), .B2(new_n795), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1212), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n792), .A2(new_n1168), .B1(new_n1069), .B2(new_n782), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT114), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n810), .A2(G128), .B1(new_n801), .B2(new_n1172), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n854), .B2(new_n793), .C1(new_n849), .C2(new_n795), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1224), .B1(new_n777), .B2(new_n774), .C1(new_n1229), .C2(KEYINPUT59), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1211), .B1(new_n1232), .B2(new_n764), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1209), .A2(new_n754), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1160), .A2(new_n1145), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT57), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n702), .B1(new_n1235), .B2(KEYINPUT57), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(G375));
  INV_X1    g1038(.A(KEYINPUT115), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1143), .A2(new_n832), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n946), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1138), .B1(new_n748), .B2(new_n915), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1240), .A2(new_n1122), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1239), .B1(new_n1244), .B2(new_n753), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1159), .A2(KEYINPUT115), .A3(new_n754), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n975), .A2(G294), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n810), .A2(G283), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n845), .A2(new_n776), .B1(new_n773), .B2(new_n205), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1067), .A2(new_n248), .A3(new_n1249), .A4(new_n980), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G107), .A2(new_n843), .B1(new_n808), .B2(G116), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G128), .A2(new_n785), .B1(new_n801), .B2(G159), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n202), .B2(new_n782), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n401), .B1(new_n799), .B2(G58), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(KEYINPUT116), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G150), .A2(new_n843), .B1(new_n808), .B2(new_n1172), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(KEYINPUT116), .A2(new_n1255), .B1(new_n810), .B2(G137), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n792), .A2(new_n854), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1252), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n764), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1263), .B(new_n755), .C1(G68), .C2(new_n838), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n946), .B2(new_n766), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1245), .A2(new_n1246), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1022), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n952), .A2(new_n1144), .A3(new_n668), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1156), .A2(new_n1269), .A3(new_n1158), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1153), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(G381));
  OR2_X1    g1073(.A1(G375), .A2(KEYINPUT117), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G375), .A2(KEYINPUT117), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1161), .A2(new_n1162), .A3(new_n1185), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n996), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1040), .B1(new_n1050), .B2(new_n754), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT108), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1278), .B1(new_n1281), .B2(new_n1051), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1277), .A2(new_n1282), .A3(new_n1272), .A4(new_n1283), .ZN(G407));
  NAND2_X1  g1084(.A1(new_n674), .A2(G213), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G407), .A2(G213), .A3(new_n1287), .ZN(G409));
  OAI21_X1  g1088(.A(new_n1145), .B1(new_n1142), .B2(new_n1153), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1209), .A3(new_n1268), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT118), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1210), .A2(new_n1233), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT119), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1201), .A2(new_n1192), .A3(new_n1202), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1206), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1203), .A2(new_n1208), .A3(KEYINPUT119), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n754), .A3(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1289), .A2(new_n1209), .A3(KEYINPUT118), .A4(new_n1268), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1292), .A2(new_n1293), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1276), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1234), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1286), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G384), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1269), .A4(new_n1158), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1153), .A2(new_n1306), .A3(new_n702), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT60), .B1(new_n1244), .B2(new_n1269), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1305), .B1(new_n1309), .B2(new_n1267), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1270), .A2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1312), .A2(new_n702), .A3(new_n1153), .A4(new_n1306), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1159), .A2(new_n754), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1265), .B1(new_n1314), .B2(new_n1239), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1313), .A2(new_n1315), .A3(G384), .A4(new_n1246), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1304), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT63), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT124), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1118), .B1(new_n1119), .B2(new_n753), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(G387), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n996), .B(G390), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT123), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT124), .B1(new_n1282), .B2(G390), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1282), .A2(KEYINPUT123), .A3(G390), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1325), .A2(new_n1328), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(G393), .B(G396), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT125), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1332), .B1(new_n1282), .B2(G390), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1326), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(new_n1324), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1339), .A2(KEYINPUT125), .A3(new_n1332), .A4(new_n1326), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT61), .B1(new_n1334), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT120), .ZN(new_n1344));
  INV_X1    g1144(.A(G2897), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1285), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1346), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1310), .A2(new_n1316), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT121), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1310), .A2(KEYINPUT121), .A3(new_n1316), .A4(new_n1347), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1285), .A2(new_n1345), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1317), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT122), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1304), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  AOI22_X1  g1157(.A1(new_n1350), .A2(new_n1351), .B1(new_n1317), .B2(new_n1353), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(KEYINPUT122), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1343), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1321), .B(new_n1342), .C1(new_n1360), .C2(new_n1320), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1334), .A2(new_n1362), .A3(new_n1341), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1362), .B1(new_n1334), .B2(new_n1341), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT61), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1366), .B1(new_n1355), .B2(new_n1304), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT62), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1319), .A2(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1304), .A2(KEYINPUT62), .A3(new_n1318), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1367), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1365), .B1(new_n1371), .B2(KEYINPUT126), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1304), .ZN(new_n1373));
  AOI21_X1  g1173(.A(KEYINPUT61), .B1(new_n1373), .B2(new_n1358), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1370), .ZN(new_n1375));
  AOI21_X1  g1175(.A(KEYINPUT62), .B1(new_n1304), .B2(new_n1318), .ZN(new_n1376));
  OAI211_X1 g1176(.A(new_n1374), .B(KEYINPUT126), .C1(new_n1375), .C2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1361), .B1(new_n1372), .B2(new_n1378), .ZN(G405));
  NAND2_X1  g1179(.A1(G375), .A2(new_n1276), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1380), .A2(new_n1303), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1318), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1365), .B(new_n1382), .ZN(G402));
endmodule


