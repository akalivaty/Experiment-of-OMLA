//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT1), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(G120gat), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n205), .A2(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n203), .A2(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT69), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n207), .A2(new_n210), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G113gat), .B2(G120gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(G120gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n225), .A2(KEYINPUT70), .A3(new_n207), .A4(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n210), .B1(new_n208), .B2(new_n209), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n203), .B2(G134gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n205), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n215), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G141gat), .B(G148gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n238), .C1(new_n239), .C2(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(G141gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G148gat), .ZN(new_n242));
  INV_X1    g041(.A(G148gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G141gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(new_n235), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  INV_X1    g052(.A(new_n249), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n227), .A2(new_n253), .A3(new_n254), .A4(new_n233), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n233), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(new_n219), .B2(new_n226), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n258), .B2(new_n254), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n252), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT78), .Z(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n254), .B1(new_n227), .B2(new_n233), .ZN(new_n265));
  AOI211_X1 g064(.A(new_n257), .B(new_n249), .C1(new_n219), .C2(new_n226), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT80), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(KEYINPUT5), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n262), .B1(new_n234), .B2(new_n251), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n254), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n255), .A2(KEYINPUT79), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n264), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n264), .B(KEYINPUT84), .C1(new_n271), .C2(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n264), .B(new_n287), .C1(new_n271), .C2(new_n279), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n259), .B1(KEYINPUT79), .B2(new_n255), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n274), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n272), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n268), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n287), .B1(new_n299), .B2(new_n264), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n290), .A2(new_n294), .B1(KEYINPUT6), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n303));
  AOI21_X1  g102(.A(G190gat), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT25), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT25), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n307), .B(new_n308), .C1(G183gat), .C2(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT27), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n325), .A2(new_n326), .A3(G190gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT64), .B(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n321), .A3(G183gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(KEYINPUT65), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n327), .B1(new_n334), .B2(new_n326), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(KEYINPUT66), .A3(new_n338), .A4(new_n313), .ZN(new_n339));
  NOR3_X1   g138(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n342), .A3(new_n305), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n317), .B(new_n320), .C1(new_n335), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n258), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n317), .A2(new_n320), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n333), .A2(new_n330), .A3(new_n332), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n321), .B1(new_n302), .B2(new_n303), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n326), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n327), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n234), .ZN(new_n353));
  NAND2_X1  g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n345), .A2(new_n353), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n354), .ZN(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G43gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT72), .B(G15gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT34), .B1(new_n355), .B2(KEYINPUT73), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n356), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n359), .B(new_n354), .C1(new_n357), .C2(new_n364), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n366), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n366), .A2(new_n372), .B1(new_n370), .B2(new_n371), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n380));
  AND2_X1   g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  OR2_X1    g180(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(G197gat), .A2(G204gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  NOR2_X1   g188(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G197gat), .B(G204gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT75), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n388), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n393), .A3(new_n394), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n379), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n394), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n402), .B2(new_n380), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT76), .B1(new_n403), .B2(new_n395), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n378), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n254), .B1(new_n405), .B2(new_n250), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n254), .B2(new_n250), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n408), .A2(new_n401), .A3(new_n404), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n377), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n402), .B(new_n399), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n250), .B1(new_n411), .B2(new_n407), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n377), .B1(new_n412), .B2(new_n249), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n401), .A2(new_n404), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(new_n408), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(G22gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT31), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G50gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n410), .A2(new_n419), .A3(new_n416), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n419), .B1(new_n410), .B2(new_n416), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n376), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n344), .B2(new_n378), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n352), .A2(new_n433), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n435), .A2(new_n436), .A3(new_n414), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n352), .B2(new_n407), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n344), .A2(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n415), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n432), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n407), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n344), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n414), .B1(new_n443), .B2(new_n436), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n439), .B(new_n415), .C1(new_n445), .C2(new_n434), .ZN(new_n446));
  INV_X1    g245(.A(new_n432), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(new_n440), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT35), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT82), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OR3_X1    g257(.A1(new_n301), .A2(new_n429), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n280), .A2(new_n288), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n292), .A3(new_n291), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n280), .A2(KEYINPUT6), .A3(new_n288), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(new_n452), .B2(new_n449), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n366), .A2(new_n372), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n370), .A2(new_n371), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND4_X1   g266(.A1(new_n424), .A2(new_n428), .A3(new_n373), .A4(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n460), .B(new_n456), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n428), .A2(new_n424), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n463), .B1(new_n293), .B2(new_n300), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n453), .A4(new_n376), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT86), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n459), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n455), .A2(new_n457), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n265), .A2(new_n266), .A3(new_n262), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n477), .B(new_n478), .C1(new_n260), .C2(new_n262), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n260), .A2(new_n477), .A3(new_n262), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n287), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n482), .B2(KEYINPUT40), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT83), .B(new_n484), .C1(new_n479), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n290), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n470), .B1(new_n475), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n447), .B1(new_n450), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n489), .B2(new_n450), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT38), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n290), .A2(new_n294), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n438), .A2(new_n439), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n489), .B1(new_n495), .B2(new_n415), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n439), .B(new_n414), .C1(new_n445), .C2(new_n434), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT38), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n490), .A2(new_n498), .B1(new_n450), .B2(new_n447), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n463), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n493), .B1(new_n500), .B2(KEYINPUT85), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n301), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n488), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n376), .B(KEYINPUT36), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n464), .B2(new_n470), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n474), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT91), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n508), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT7), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(G92gat), .ZN(new_n515));
  INV_X1    g314(.A(G85gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n515), .A2(new_n516), .B1(KEYINPUT8), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G99gat), .B(G106gat), .Z(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G57gat), .B(G64gat), .Z(new_n524));
  INV_X1    g323(.A(G71gat), .ZN(new_n525));
  INV_X1    g324(.A(G78gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(KEYINPUT9), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G71gat), .B(G78gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT10), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n521), .A2(new_n530), .A3(new_n522), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT94), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n532), .A2(new_n537), .A3(new_n533), .A4(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT10), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n542), .B1(new_n532), .B2(new_n534), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(KEYINPUT95), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n543), .B(new_n548), .C1(KEYINPUT95), .C2(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(new_n542), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n535), .A2(KEYINPUT94), .B1(KEYINPUT10), .B2(new_n539), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n538), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n552), .B2(new_n547), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n553), .A2(KEYINPUT96), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(KEYINPUT96), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT13), .Z(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n561));
  AOI211_X1 g360(.A(new_n560), .B(new_n561), .C1(G29gat), .C2(G36gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT14), .ZN(new_n563));
  INV_X1    g362(.A(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(KEYINPUT88), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n567), .A2(KEYINPUT87), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n567), .B2(KEYINPUT87), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n572), .A2(new_n573), .B1(new_n564), .B2(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n561), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(G1gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(G1gat), .B2(new_n578), .ZN(new_n581));
  INV_X1    g380(.A(G8gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(KEYINPUT89), .A3(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT89), .B1(new_n577), .B2(new_n583), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n558), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n571), .A2(KEYINPUT17), .A3(new_n575), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n592), .A3(new_n557), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n584), .A2(new_n592), .A3(KEYINPUT18), .A4(new_n557), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G197gat), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT11), .B(G169gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n595), .A3(new_n596), .A4(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n556), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n507), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n392), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n523), .A3(new_n591), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n576), .A2(new_n521), .A3(new_n522), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n622), .B(new_n613), .C1(new_n617), .C2(new_n618), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n621), .A2(new_n330), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n330), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G190gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n330), .A3(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n611), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n583), .B1(new_n633), .B2(new_n531), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n530), .B(KEYINPUT21), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n635), .B2(new_n583), .ZN(new_n636));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G127gat), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n641), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n632), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n471), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT97), .B(G1gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  NOR2_X1   g453(.A1(new_n648), .A2(new_n475), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n655), .B2(new_n582), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  MUX2_X1   g457(.A(KEYINPUT42), .B(new_n656), .S(new_n658), .Z(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n648), .A2(new_n660), .A3(new_n505), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n376), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n660), .B2(new_n662), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n470), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n631), .A2(new_n645), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n609), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n564), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n609), .A2(KEYINPUT100), .A3(new_n668), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n674));
  AND3_X1   g473(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n671), .B2(new_n673), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n631), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n503), .A3(new_n492), .ZN(new_n683));
  INV_X1    g482(.A(new_n488), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n506), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n301), .A2(new_n429), .A3(new_n458), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n460), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n472), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n681), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n646), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n464), .B2(new_n470), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n471), .A2(new_n453), .ZN(new_n695));
  INV_X1    g494(.A(new_n470), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT101), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n697), .A3(new_n505), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n474), .B1(new_n504), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n699), .B2(new_n632), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n679), .B1(new_n701), .B2(new_n608), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n683), .B2(new_n684), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n632), .B1(new_n703), .B2(new_n690), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n680), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n645), .B1(new_n507), .B2(new_n681), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n679), .A2(new_n705), .A3(new_n608), .A4(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n678), .B(new_n650), .C1(new_n702), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G29gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n701), .A2(new_n679), .A3(new_n608), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n608), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n678), .B1(new_n713), .B2(new_n650), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n677), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT104), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(new_n677), .C1(new_n709), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1328gat));
  NOR3_X1   g518(.A1(new_n669), .A2(G36gat), .A3(new_n475), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n475), .B1(new_n710), .B2(new_n712), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n565), .ZN(G1329gat));
  INV_X1    g522(.A(new_n376), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n669), .A2(G43gat), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n711), .B2(new_n505), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n505), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n725), .B1(new_n730), .B2(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n731), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n696), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n609), .A2(new_n668), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n470), .B1(new_n710), .B2(new_n712), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n733), .B(new_n737), .C1(new_n738), .C2(new_n734), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n740));
  OAI21_X1  g539(.A(G50gat), .B1(new_n711), .B2(new_n470), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT48), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n740), .B1(new_n739), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  AND2_X1   g545(.A1(new_n699), .A2(new_n607), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n647), .A3(new_n556), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n471), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT107), .B(G57gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT108), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n749), .B(new_n751), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n748), .A2(new_n475), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  AND2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n753), .B2(new_n754), .ZN(G1333gat));
  OR3_X1    g556(.A1(new_n748), .A2(new_n525), .A3(new_n505), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n525), .B1(new_n748), .B2(new_n724), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT50), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1334gat));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n647), .A3(new_n556), .A4(new_n696), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g566(.A1(new_n747), .A2(new_n668), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n556), .A2(new_n516), .A3(new_n650), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(new_n556), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n692), .A2(new_n700), .A3(new_n606), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n650), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n775), .A2(new_n777), .B1(new_n516), .B2(new_n780), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  INV_X1    g581(.A(new_n475), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n515), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n778), .A2(G92gat), .A3(new_n475), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n782), .B(new_n786), .C1(new_n775), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n784), .B2(new_n785), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n768), .B(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n787), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n790), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n796), .B2(new_n782), .ZN(G1337gat));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n729), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G99gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n778), .A2(new_n724), .A3(G99gat), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT114), .Z(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n775), .B2(new_n801), .ZN(G1338gat));
  NAND2_X1  g601(.A1(new_n779), .A2(new_n696), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n778), .A2(G106gat), .A3(new_n470), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n794), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n773), .B2(new_n774), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n803), .B2(G106gat), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(G1339gat));
  OAI21_X1  g613(.A(KEYINPUT117), .B1(new_n541), .B2(new_n542), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n551), .A2(new_n816), .A3(new_n550), .A4(new_n538), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n543), .A4(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n546), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n552), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n549), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n821), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n606), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n586), .A2(new_n558), .A3(new_n587), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n557), .B1(new_n584), .B2(new_n592), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n601), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n556), .A2(new_n605), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n632), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n823), .A2(new_n826), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n605), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n605), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n626), .A2(new_n630), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n646), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n632), .A2(new_n646), .A3(new_n606), .A4(new_n556), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n429), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n783), .A2(new_n471), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n606), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G113gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n224), .B2(new_n846), .ZN(G1340gat));
  NAND2_X1  g647(.A1(new_n556), .A2(new_n209), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT119), .Z(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n845), .A2(new_n556), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n209), .ZN(G1341gat));
  NAND2_X1  g652(.A1(new_n845), .A2(new_n645), .ZN(new_n854));
  XOR2_X1   g653(.A(KEYINPUT120), .B(G127gat), .Z(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1342gat));
  AND2_X1   g655(.A1(new_n845), .A2(new_n632), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n205), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n205), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(KEYINPUT56), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(KEYINPUT56), .B2(new_n859), .ZN(G1343gat));
  AND3_X1   g660(.A1(new_n626), .A2(new_n630), .A3(new_n837), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n823), .A3(new_n826), .A4(new_n835), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n553), .B(KEYINPUT96), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n834), .B1(new_n864), .B2(new_n549), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT121), .B1(new_n824), .B2(new_n825), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(KEYINPUT55), .C1(new_n818), .C2(new_n821), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n606), .A2(new_n822), .A3(new_n549), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n871), .B2(new_n632), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n841), .B1(new_n872), .B2(new_n646), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n470), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n840), .A2(new_n842), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n696), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n505), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n874), .A2(new_n606), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G141gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n607), .A2(G141gat), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n875), .A2(new_n696), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT123), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n888), .B(new_n885), .C1(new_n880), .C2(G141gat), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n470), .B1(new_n840), .B2(new_n842), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n879), .A4(new_n882), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(G141gat), .B2(new_n880), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n887), .A2(new_n889), .B1(new_n895), .B2(new_n884), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT124), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  OAI221_X1 g697(.A(new_n898), .B1(new_n895), .B2(new_n884), .C1(new_n887), .C2(new_n889), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(new_n892), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n878), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n243), .A3(new_n556), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n874), .A2(new_n877), .A3(new_n879), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n243), .C1(new_n905), .C2(new_n556), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n873), .A2(new_n470), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n556), .A3(new_n879), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n906), .B2(new_n912), .ZN(G1345gat));
  AOI21_X1  g712(.A(G155gat), .B1(new_n902), .B2(new_n645), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n646), .A2(new_n236), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n905), .B2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n904), .B2(new_n631), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n237), .A3(new_n632), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n475), .A2(new_n429), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(new_n650), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n875), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G169gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n606), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n475), .A2(new_n650), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n843), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n606), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n926), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n925), .B2(new_n556), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n556), .A2(G176gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n929), .B2(new_n933), .ZN(G1349gat));
  AOI21_X1  g733(.A(new_n328), .B1(new_n929), .B2(new_n645), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n924), .A2(new_n646), .A3(new_n325), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g737(.A(new_n330), .B1(new_n929), .B2(new_n632), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT61), .Z(new_n940));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n330), .A3(new_n632), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1351gat));
  NAND2_X1  g741(.A1(new_n928), .A2(new_n505), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n901), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g743(.A(KEYINPUT126), .B(G197gat), .Z(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n606), .A3(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n910), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n607), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n945), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n951), .A3(new_n556), .ZN(new_n952));
  XOR2_X1   g751(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n910), .A2(new_n556), .A3(new_n947), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n951), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n944), .A2(new_n391), .A3(new_n645), .ZN(new_n957));
  INV_X1    g756(.A(new_n948), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n645), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n944), .B2(new_n632), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n631), .A2(new_n392), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n958), .B2(new_n964), .ZN(G1355gat));
endmodule


