//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205));
  INV_X1    g004(.A(G85gat), .ZN(new_n206));
  INV_X1    g005(.A(G92gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(KEYINPUT8), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n206), .A2(new_n207), .B1(new_n209), .B2(KEYINPUT96), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n211), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G99gat), .B(G106gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT97), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n208), .A2(new_n214), .A3(new_n210), .A4(new_n212), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G71gat), .ZN(new_n223));
  INV_X1    g022(.A(G78gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(KEYINPUT9), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT94), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT93), .ZN(new_n230));
  INV_X1    g029(.A(G64gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(G57gat), .ZN(new_n232));
  INV_X1    g031(.A(G57gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT93), .B1(new_n233), .B2(G64gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(G64gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n232), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n230), .B1(new_n231), .B2(G57gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(G57gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n229), .B1(new_n240), .B2(new_n232), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n228), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(G64gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR3_X1   g046(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n248));
  NOR4_X1   g047(.A1(new_n245), .A2(new_n225), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT95), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT94), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n227), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n254), .A2(new_n255), .A3(new_n249), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n222), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT100), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n242), .A2(new_n250), .A3(new_n218), .A4(new_n216), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n222), .B(KEYINPUT100), .C1(new_n251), .C2(new_n256), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n251), .A2(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n204), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n204), .ZN(new_n269));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G204gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n267), .B2(new_n269), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n264), .A2(KEYINPUT21), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n264), .A2(KEYINPUT21), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT16), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(G1gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n287), .B(new_n288), .C1(G1gat), .C2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(G8gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n281), .B(G127gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n298));
  XNOR2_X1  g097(.A(G155gat), .B(G183gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(G211gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n300), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n293), .A2(new_n296), .A3(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G43gat), .B(G50gat), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT15), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(G29gat), .A2(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT14), .ZN(new_n314));
  NAND2_X1  g113(.A1(G29gat), .A2(G36gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n315), .B(KEYINPUT84), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n320), .A2(new_n323), .B1(new_n311), .B2(new_n310), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n312), .A2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(KEYINPUT86), .A3(new_n325), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n319), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n330), .A2(KEYINPUT87), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n324), .A2(KEYINPUT86), .A3(new_n325), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT86), .B1(new_n324), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n318), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT17), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n222), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G232gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n338), .A2(KEYINPUT98), .B1(KEYINPUT41), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n331), .B1(new_n330), .B2(KEYINPUT87), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT17), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT98), .B(new_n221), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G190gat), .B(G218gat), .Z(new_n346));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n222), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n341), .A2(new_n345), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT99), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n345), .A3(new_n348), .ZN(new_n351));
  INV_X1    g150(.A(new_n346), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n340), .A2(KEYINPUT41), .ZN(new_n354));
  XNOR2_X1  g153(.A(G134gat), .B(G162gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n353), .A3(new_n349), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n356), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n309), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT27), .B(G183gat), .Z(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT64), .B(G190gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366));
  OR4_X1    g165(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(G169gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n271), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT66), .B1(new_n369), .B2(KEYINPUT26), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(KEYINPUT26), .ZN(new_n371));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n367), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT65), .B(KEYINPUT28), .C1(new_n362), .C2(new_n363), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n365), .A2(new_n366), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OR3_X1    g174(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n376), .A2(new_n377), .B1(G169gat), .B2(G176gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n363), .A2(G183gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n366), .B(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT25), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n384));
  NOR2_X1   g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n378), .B(new_n384), .C1(new_n381), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n375), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT67), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n388), .A2(new_n282), .A3(G134gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT1), .ZN(new_n393));
  MUX2_X1   g192(.A(new_n391), .B(new_n390), .S(new_n393), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n383), .A2(new_n386), .ZN(new_n398));
  INV_X1    g197(.A(new_n394), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n375), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n394), .A3(KEYINPUT68), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT32), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  XNOR2_X1  g205(.A(G15gat), .B(G43gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(G71gat), .ZN(new_n408));
  INV_X1    g207(.A(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  OAI221_X1 g211(.A(KEYINPUT32), .B1(new_n405), .B2(new_n412), .C1(new_n402), .C2(new_n403), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n397), .A2(new_n400), .A3(new_n403), .A4(new_n401), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT34), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n414), .A2(new_n416), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(KEYINPUT71), .A3(new_n416), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G57gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G85gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427));
  OR2_X1    g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(KEYINPUT2), .ZN(new_n429));
  XOR2_X1   g228(.A(G141gat), .B(G148gat), .Z(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n427), .A3(new_n428), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT4), .B1(new_n437), .B2(new_n394), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n431), .B(KEYINPUT77), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n399), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(KEYINPUT3), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n433), .A2(new_n447), .A3(new_n436), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n394), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(new_n399), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n394), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n445), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n399), .B1(new_n441), .B2(new_n447), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n446), .A2(new_n456), .B1(new_n438), .B2(new_n443), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n445), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n426), .B(new_n452), .C1(new_n458), .C2(new_n451), .ZN(new_n459));
  INV_X1    g258(.A(new_n426), .ZN(new_n460));
  INV_X1    g259(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n451), .B1(new_n450), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT5), .B1(new_n457), .B2(new_n445), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n426), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(new_n231), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(new_n207), .ZN(new_n472));
  XOR2_X1   g271(.A(G211gat), .B(G218gat), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G211gat), .A2(G218gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT22), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G197gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n273), .ZN(new_n479));
  NOR2_X1   g278(.A1(G197gat), .A2(G204gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n474), .A2(KEYINPUT72), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n474), .B1(new_n481), .B2(KEYINPUT72), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G226gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(new_n203), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n398), .A2(new_n489), .A3(new_n375), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n387), .A2(KEYINPUT73), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n487), .A2(KEYINPUT29), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n398), .B2(new_n375), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n485), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n398), .A2(new_n487), .A3(new_n375), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n490), .A2(new_n491), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n484), .B(new_n497), .C1(new_n498), .C2(new_n494), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n472), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OR3_X1    g299(.A1(new_n500), .A2(KEYINPUT76), .A3(KEYINPUT30), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n472), .B(KEYINPUT75), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n496), .A2(KEYINPUT74), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT74), .B1(new_n496), .B2(new_n499), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT30), .B1(new_n500), .B2(KEYINPUT76), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n469), .A2(new_n507), .A3(KEYINPUT35), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(G22gat), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n437), .A2(new_n484), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n446), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n448), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n485), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(KEYINPUT80), .A3(new_n446), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G228gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n203), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n481), .B1(KEYINPUT78), .B2(new_n473), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n473), .A2(KEYINPUT78), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n512), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n447), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n437), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(new_n518), .C1(new_n521), .C2(new_n203), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n523), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n523), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n511), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n533), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n510), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n422), .A2(new_n508), .A3(KEYINPUT82), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n419), .A2(new_n543), .A3(new_n420), .A4(new_n421), .ZN(new_n546));
  INV_X1    g345(.A(new_n507), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n466), .A2(new_n468), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n469), .A2(new_n507), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n416), .A2(KEYINPUT69), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n414), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n411), .A2(KEYINPUT69), .A3(new_n416), .A4(new_n413), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n555), .A2(new_n556), .B1(new_n538), .B2(new_n542), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n548), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n564));
  INV_X1    g363(.A(new_n553), .ZN(new_n565));
  INV_X1    g364(.A(new_n543), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n562), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT37), .B1(new_n496), .B2(new_n499), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT81), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n492), .A2(new_n495), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n484), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n497), .B1(new_n498), .B2(new_n494), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n485), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT38), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(new_n502), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT37), .B1(new_n503), .B2(new_n504), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n569), .A2(new_n472), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n500), .A2(KEYINPUT38), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n469), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n444), .A2(new_n449), .ZN(new_n581));
  INV_X1    g380(.A(new_n445), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n453), .A2(new_n454), .A3(new_n445), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(KEYINPUT39), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n585), .B(new_n460), .C1(KEYINPUT39), .C2(new_n583), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT40), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n459), .A3(new_n507), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(new_n543), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n552), .A2(new_n559), .B1(new_n567), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n291), .B1(new_n332), .B2(new_n337), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n330), .A2(new_n291), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT89), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n330), .B(new_n291), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(KEYINPUT90), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n592), .A2(KEYINPUT18), .A3(new_n593), .A4(new_n595), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n598), .A2(new_n612), .A3(new_n602), .A4(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n591), .A2(KEYINPUT91), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n611), .A2(new_n613), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n590), .B2(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n280), .B(new_n361), .C1(new_n615), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n469), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT102), .B(G1gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(G1324gat));
  NAND2_X1  g421(.A1(new_n286), .A2(new_n290), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n619), .A2(new_n507), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n615), .A2(new_n618), .ZN(new_n629));
  INV_X1    g428(.A(new_n361), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n279), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(G8gat), .B1(new_n631), .B2(new_n547), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT103), .B1(new_n633), .B2(new_n625), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n625), .A2(new_n627), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(G1325gat));
  NAND2_X1  g435(.A1(new_n562), .A2(new_n564), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n619), .A2(G15gat), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(G15gat), .B1(new_n619), .B2(new_n422), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(G1326gat));
  NAND2_X1  g443(.A1(new_n619), .A2(new_n566), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n309), .A2(new_n280), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n360), .A2(new_n357), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT105), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n549), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT106), .B1(new_n552), .B2(new_n559), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  AOI211_X1 g456(.A(new_n657), .B(new_n558), .C1(new_n544), .C2(new_n551), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n567), .A2(new_n589), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n649), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n590), .A2(new_n655), .A3(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n662), .A2(new_n614), .A3(new_n648), .A4(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n665), .A2(new_n666), .A3(new_n549), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n665), .B2(new_n549), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(G29gat), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n669), .ZN(G1328gat));
  NOR3_X1   g469(.A1(new_n652), .A2(G36gat), .A3(new_n547), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT46), .ZN(new_n672));
  OAI21_X1  g471(.A(G36gat), .B1(new_n665), .B2(new_n547), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  OAI21_X1  g473(.A(G43gat), .B1(new_n665), .B2(new_n637), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT47), .B1(new_n675), .B2(KEYINPUT109), .ZN(new_n676));
  INV_X1    g475(.A(G43gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n629), .A2(new_n651), .A3(new_n677), .A4(new_n422), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n678), .B(KEYINPUT108), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n684), .B(new_n675), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n665), .B2(new_n543), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT48), .B1(new_n687), .B2(KEYINPUT111), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n543), .A2(G50gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT110), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n629), .A2(new_n651), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n687), .B(new_n691), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1331gat));
  NOR3_X1   g494(.A1(new_n660), .A2(new_n614), .A3(new_n361), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n280), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n549), .B(KEYINPUT112), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n233), .ZN(G1332gat));
  AND2_X1   g500(.A1(new_n696), .A2(new_n280), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT114), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n547), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT113), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n707), .A2(new_n708), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n708), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n706), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(G1333gat));
  NAND3_X1  g512(.A1(new_n702), .A2(G71gat), .A3(new_n638), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n223), .B1(new_n697), .B2(new_n560), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g516(.A1(new_n697), .A2(new_n543), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n224), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n309), .A2(new_n614), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n662), .A2(new_n280), .A3(new_n664), .A4(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(new_n206), .A3(new_n549), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n552), .A2(new_n559), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n657), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n567), .A2(new_n589), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n552), .A2(KEYINPUT106), .A3(new_n559), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n649), .A3(new_n720), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT51), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n727), .A2(new_n730), .A3(new_n649), .A4(new_n720), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n729), .A2(new_n469), .A3(new_n280), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n722), .B1(new_n206), .B2(new_n732), .ZN(G1336gat));
  NOR2_X1   g532(.A1(new_n547), .A2(G92gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n729), .A2(new_n280), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n721), .A2(new_n547), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n207), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT52), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n739), .B(new_n735), .C1(new_n736), .C2(new_n207), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n721), .B2(new_n637), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n729), .A2(new_n409), .A3(new_n280), .A4(new_n731), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n560), .B2(new_n743), .ZN(G1338gat));
  INV_X1    g543(.A(G106gat), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n727), .B2(new_n649), .ZN(new_n746));
  INV_X1    g545(.A(new_n720), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n746), .A2(new_n279), .A3(new_n663), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(new_n566), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n280), .A3(new_n566), .A4(new_n731), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT53), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(KEYINPUT115), .A3(new_n566), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n721), .B2(new_n543), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n755), .A3(G106gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n750), .B2(G106gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n752), .B1(new_n756), .B2(new_n758), .ZN(G1339gat));
  NOR3_X1   g558(.A1(new_n361), .A2(new_n280), .A3(new_n614), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n263), .A2(new_n265), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  INV_X1    g562(.A(new_n204), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n263), .A2(new_n204), .A3(new_n265), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT54), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n274), .B(new_n765), .C1(new_n767), .C2(new_n266), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n276), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n267), .A2(KEYINPUT54), .A3(new_n766), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n275), .B1(new_n266), .B2(new_n763), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n761), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n769), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(KEYINPUT55), .A3(new_n772), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT116), .A4(new_n276), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n599), .A2(new_n601), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n609), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n613), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n649), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(new_n279), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n778), .B2(new_n614), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(new_n649), .ZN(new_n787));
  INV_X1    g586(.A(new_n309), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n760), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n699), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n547), .ZN(new_n791));
  INV_X1    g590(.A(new_n557), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(G113gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n614), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n789), .B2(new_n566), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n617), .B1(new_n774), .B2(new_n777), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n661), .B1(new_n798), .B2(new_n785), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n309), .B1(new_n799), .B2(new_n784), .ZN(new_n800));
  OAI211_X1 g599(.A(KEYINPUT117), .B(new_n543), .C1(new_n800), .C2(new_n760), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n560), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n507), .A2(new_n549), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n614), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n795), .B1(new_n805), .B2(new_n794), .ZN(G1340gat));
  INV_X1    g605(.A(G120gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n793), .A2(new_n807), .A3(new_n280), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n804), .A2(new_n280), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1341gat));
  AOI21_X1  g609(.A(G127gat), .B1(new_n793), .B2(new_n309), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n788), .A2(new_n282), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n804), .B2(new_n812), .ZN(G1342gat));
  NAND2_X1  g612(.A1(new_n649), .A2(new_n547), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT118), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n814), .A2(KEYINPUT118), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n790), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(G134gat), .A3(new_n792), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT56), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n649), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G134gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1343gat));
  INV_X1    g621(.A(G141gat), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n768), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n614), .A2(new_n276), .A3(new_n776), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n785), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n661), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n784), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n760), .B1(new_n830), .B2(new_n788), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n831), .B2(new_n543), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n566), .C1(new_n800), .C2(new_n760), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n637), .A2(new_n803), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT119), .Z(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n832), .A2(new_n839), .A3(new_n834), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n823), .B1(new_n841), .B2(new_n614), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n638), .A2(new_n543), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n791), .A2(G141gat), .A3(new_n617), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT58), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n847));
  OAI21_X1  g646(.A(G141gat), .B1(new_n837), .B2(new_n617), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(G1344gat));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n770), .A2(new_n773), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n649), .A2(new_n852), .A3(new_n783), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n649), .B1(new_n827), .B2(new_n826), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n788), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n760), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n543), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n566), .C1(new_n800), .C2(new_n760), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n829), .A2(new_n853), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n760), .B1(new_n861), .B2(new_n788), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT122), .B(new_n833), .C1(new_n862), .C2(new_n543), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n280), .A3(new_n836), .ZN(new_n865));
  AND2_X1   g664(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n791), .A2(new_n844), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n279), .A2(G148gat), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(G148gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n841), .B2(new_n280), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g671(.A(G155gat), .B1(new_n867), .B2(new_n309), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n788), .B1(new_n838), .B2(new_n840), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g674(.A(new_n661), .B1(new_n838), .B2(new_n840), .ZN(new_n876));
  INV_X1    g675(.A(G162gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n843), .A2(new_n877), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n876), .A2(new_n877), .B1(new_n817), .B2(new_n878), .ZN(G1347gat));
  NOR4_X1   g678(.A1(new_n789), .A2(new_n469), .A3(new_n547), .A4(new_n792), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n368), .A3(new_n614), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n699), .A2(new_n507), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT123), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n802), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n614), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n885), .B2(new_n368), .ZN(G1348gat));
  AOI21_X1  g685(.A(G176gat), .B1(new_n880), .B2(new_n280), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n279), .A2(new_n271), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(G1349gat));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890));
  INV_X1    g689(.A(new_n880), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(new_n362), .A3(new_n788), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n884), .A2(new_n309), .ZN(new_n894));
  INV_X1    g693(.A(G183gat), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n890), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n884), .B2(new_n309), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n897), .B2(new_n892), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1350gat));
  NAND2_X1  g698(.A1(new_n797), .A2(new_n801), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(new_n422), .A3(new_n649), .A4(new_n883), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G190gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n905));
  INV_X1    g704(.A(new_n363), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n906), .A3(new_n649), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n880), .A2(new_n909), .A3(new_n906), .A4(new_n649), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n904), .A2(new_n914), .A3(new_n905), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n864), .A2(new_n637), .A3(new_n883), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n617), .ZN(new_n918));
  NOR4_X1   g717(.A1(new_n789), .A2(new_n844), .A3(new_n469), .A4(new_n547), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n478), .A3(new_n614), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1352gat));
  OR3_X1    g720(.A1(new_n917), .A2(KEYINPUT126), .A3(new_n279), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT126), .B1(new_n917), .B2(new_n279), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(G204gat), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(new_n273), .A3(new_n280), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT62), .Z(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n919), .A2(new_n303), .A3(new_n309), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n864), .A2(new_n637), .A3(new_n309), .A4(new_n883), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1354gat));
  INV_X1    g731(.A(G218gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n933), .A3(new_n649), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n661), .B1(new_n917), .B2(KEYINPUT127), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n864), .A2(new_n936), .A3(new_n637), .A4(new_n883), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n938), .B2(new_n933), .ZN(G1355gat));
endmodule


