//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(G137), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n462), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(KEYINPUT71), .B(new_n462), .C1(new_n469), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n471), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n481), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n481), .B2(new_n466), .ZN(new_n483));
  OAI21_X1  g058(.A(G125), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(G113), .A2(G2104), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n480), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n477), .A2(new_n488), .ZN(G160));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n480), .C2(G112), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT72), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n469), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n469), .A2(new_n480), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n468), .A3(new_n466), .A4(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n470), .A2(G138), .A3(new_n471), .ZN(new_n503));
  XOR2_X1   g078(.A(KEYINPUT73), .B(KEYINPUT4), .Z(new_n504));
  OAI211_X1 g079(.A(new_n503), .B(new_n504), .C1(new_n482), .C2(new_n483), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n470), .A2(G138), .A3(new_n471), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n469), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(G164));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n510), .B2(new_n509), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n512), .A2(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n519), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NOR2_X1   g099(.A1(new_n509), .A2(new_n510), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(G51), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(new_n516), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n512), .A2(new_n538), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n521), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  NAND3_X1  g118(.A1(new_n511), .A2(G43), .A3(G543), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  AOI22_X1  g129(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n521), .B1(new_n517), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  AND2_X1   g138(.A1(new_n514), .A2(new_n515), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n525), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n527), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT74), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n514), .B2(new_n515), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT75), .B(G651), .C1(new_n571), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n565), .A2(G86), .B1(G48), .B2(new_n527), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n512), .A2(new_n583), .B1(new_n517), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n576), .B2(new_n577), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n582), .A2(new_n587), .ZN(G305));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n512), .A2(new_n589), .B1(new_n517), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n521), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n517), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT77), .B(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n564), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n527), .B2(G54), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(G868), .B2(new_n606), .ZN(G284));
  OAI21_X1  g182(.A(new_n596), .B1(G868), .B2(new_n606), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n561), .B2(G868), .ZN(G280));
  XOR2_X1   g185(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(G148));
  NOR2_X1   g188(.A1(new_n549), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n612), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n464), .A2(G2104), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n481), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n624), .A2(G2104), .A3(new_n461), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT82), .Z(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(new_n480), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n492), .B2(G135), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n494), .A2(new_n638), .A3(G123), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n638), .B1(new_n494), .B2(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  INV_X1    g218(.A(new_n642), .ZN(new_n644));
  INV_X1    g219(.A(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n629), .A2(new_n630), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n632), .A2(new_n643), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n652), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n630), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n645), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n683), .B(new_n686), .C1(new_n678), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n698), .A2(G6), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G305), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n707), .A2(new_n711), .A3(new_n715), .A4(new_n712), .ZN(new_n716));
  NOR2_X1   g291(.A1(G25), .A2(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n492), .A2(G131), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G107), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n634), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n494), .B2(G119), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n717), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n698), .A2(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n594), .B2(new_n698), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1986), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n714), .A2(new_n716), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n714), .A2(new_n738), .A3(new_n716), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n698), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G286), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n549), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G16), .B2(G19), .ZN(new_n753));
  INV_X1    g328(.A(G1341), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n750), .B(new_n755), .C1(G29), .C2(new_n644), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n698), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n606), .B2(new_n698), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT87), .B(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n753), .A2(new_n754), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n698), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G1961), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(G1961), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n756), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n768));
  NAND2_X1  g343(.A1(G162), .A2(G29), .ZN(new_n769));
  OR2_X1    g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n768), .A3(new_n770), .ZN(new_n773));
  AOI21_X1  g348(.A(G2090), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n773), .ZN(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n775), .A2(new_n776), .A3(new_n771), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n698), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NOR2_X1   g356(.A1(G27), .A2(G29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G164), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT93), .B(G2078), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n767), .A2(new_n774), .A3(new_n777), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n492), .A2(G141), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n791));
  AND3_X1   g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G129), .B2(new_n494), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G32), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT27), .B(G1996), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT24), .ZN(new_n803));
  INV_X1    g378(.A(G34), .ZN(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n803), .B2(new_n804), .ZN(new_n806));
  INV_X1    g381(.A(G29), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(G160), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G2084), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT88), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n798), .A2(new_n800), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n480), .C2(G116), .ZN(new_n814));
  INV_X1    g389(.A(new_n494), .ZN(new_n815));
  INV_X1    g390(.A(G128), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n492), .A2(G140), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n807), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n807), .A2(G33), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n624), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n480), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n492), .A2(G139), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT25), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n807), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2072), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n808), .A2(G2084), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n810), .A2(new_n823), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n787), .A2(new_n802), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n740), .A2(new_n835), .ZN(G150));
  XNOR2_X1  g411(.A(G150), .B(KEYINPUT94), .ZN(G311));
  AOI22_X1  g412(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n521), .ZN(new_n839));
  OAI211_X1 g414(.A(G55), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n517), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n606), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT95), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n549), .A2(new_n843), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n544), .B1(new_n517), .B2(new_n545), .C1(new_n547), .C2(new_n521), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n840), .B1(new_n517), .B2(new_n841), .C1(new_n838), .C2(new_n521), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n844), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n846), .B1(new_n856), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n642), .B(G160), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G162), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n797), .A2(G164), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n505), .A2(new_n507), .ZN(new_n864));
  INV_X1    g439(.A(new_n502), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n790), .A2(new_n796), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT96), .B1(new_n817), .B2(new_n818), .ZN(new_n869));
  OR3_X1    g444(.A1(new_n817), .A2(KEYINPUT96), .A3(new_n818), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n869), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n863), .A2(new_n872), .A3(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n830), .B2(KEYINPUT97), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n875), .B2(new_n830), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n878), .A3(new_n873), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n725), .B(new_n627), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n494), .A2(G130), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT99), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(KEYINPUT99), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n492), .A2(G142), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n480), .A2(G118), .ZN(new_n887));
  OAI221_X1 g462(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n887), .C2(KEYINPUT100), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(KEYINPUT100), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n725), .A2(new_n627), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n725), .A2(new_n627), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(KEYINPUT101), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n862), .B1(new_n880), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n880), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n894), .A2(KEYINPUT101), .A3(new_n897), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT101), .B1(new_n894), .B2(new_n897), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n877), .A2(new_n879), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT102), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n861), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n913));
  INV_X1    g488(.A(new_n898), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n860), .B1(new_n880), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n912), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT102), .B1(new_n908), .B2(new_n909), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n908), .A2(new_n909), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n860), .B1(new_n923), .B2(new_n910), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n915), .B2(new_n916), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT40), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n920), .A2(new_n926), .ZN(G395));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n843), .B2(G868), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n615), .B(new_n854), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n601), .A2(new_n605), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT103), .B1(new_n930), .B2(new_n561), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n606), .A2(G299), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(KEYINPUT103), .A3(new_n561), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT41), .B1(new_n938), .B2(new_n931), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n932), .A2(new_n940), .A3(new_n933), .A4(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n929), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n582), .A2(new_n587), .A3(new_n594), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G303), .B(G288), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n580), .A2(new_n581), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n948));
  AOI21_X1  g523(.A(G290), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n946), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n944), .B2(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n957));
  NAND3_X1  g532(.A1(new_n937), .A2(new_n954), .A3(new_n942), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G868), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  MUX2_X1   g537(.A(new_n928), .B(KEYINPUT105), .S(new_n962), .Z(G295));
  MUX2_X1   g538(.A(new_n928), .B(KEYINPUT105), .S(new_n962), .Z(G331));
  AND3_X1   g539(.A1(new_n850), .A2(new_n853), .A3(G301), .ZN(new_n965));
  AOI21_X1  g540(.A(G301), .B1(new_n850), .B2(new_n853), .ZN(new_n966));
  OAI21_X1  g541(.A(G286), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n549), .A2(new_n843), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n851), .A2(new_n852), .ZN(new_n969));
  OAI21_X1  g544(.A(G171), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n850), .A2(new_n853), .A3(G301), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(G168), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n939), .A2(new_n941), .A3(new_n967), .A4(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n965), .A2(new_n966), .A3(G286), .ZN(new_n974));
  AOI21_X1  g549(.A(G168), .B1(new_n970), .B2(new_n971), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n935), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n954), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(KEYINPUT106), .A3(new_n918), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n973), .A2(new_n976), .B1(new_n951), .B2(new_n953), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(G37), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n977), .B2(new_n954), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(G37), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n955), .A2(new_n976), .A3(new_n973), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI221_X1 g563(.A(KEYINPUT44), .B1(new_n983), .B2(new_n985), .C1(new_n984), .C2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n979), .A2(new_n982), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n985), .A2(G37), .A3(new_n981), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT107), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n990), .B2(KEYINPUT43), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n989), .B1(new_n996), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(G125), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n622), .B2(new_n623), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n634), .B1(new_n1004), .B2(new_n486), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(G40), .A3(new_n475), .A4(new_n476), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n819), .B(new_n821), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(G1996), .B2(new_n797), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G1996), .B2(new_n797), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n725), .B(new_n729), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1007), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n594), .B(G1986), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n866), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n1006), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n580), .A2(G1981), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n579), .B2(new_n574), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n586), .B2(new_n1025), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT49), .B1(new_n1028), .B2(KEYINPUT114), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n1021), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n703), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1021), .B1(new_n1032), .B2(new_n1024), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n703), .A2(G1976), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1021), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1021), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n1038), .A3(new_n1030), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G40), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n477), .A2(new_n488), .A3(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n468), .A2(new_n466), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n503), .A2(new_n1043), .A3(new_n465), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n506), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(KEYINPUT4), .B1(new_n624), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT45), .B(new_n1017), .C1(new_n1047), .C2(new_n502), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1048), .A3(new_n1002), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT109), .B(G1971), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n866), .A2(new_n1017), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1042), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT112), .B1(new_n1056), .B2(G2090), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G164), .A2(G1384), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1006), .B1(new_n1058), .B2(new_n1053), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n776), .A4(new_n1055), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1049), .A2(new_n1062), .A3(new_n1050), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1052), .A2(new_n1057), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1033), .B1(new_n1040), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1039), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1056), .A2(G2084), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT45), .B1(new_n866), .B2(new_n1017), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1006), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1042), .A2(KEYINPUT116), .A3(new_n1002), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1048), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1077), .B2(new_n749), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(new_n1020), .A3(G286), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1064), .A2(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1067), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1071), .A2(KEYINPUT63), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n1083));
  NOR2_X1   g658(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1083), .B(new_n1084), .C1(new_n1047), .C2(new_n502), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1053), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(G164), .B2(G1384), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1084), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(G164), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1042), .A2(new_n1085), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(G2090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1067), .B1(new_n1092), .B2(new_n1020), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(new_n1079), .A3(new_n1069), .A4(new_n1039), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1070), .B1(new_n1082), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(G299), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n561), .A2(KEYINPUT117), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1042), .A2(new_n1048), .A3(new_n1002), .A4(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1099), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1056), .A2(new_n759), .B1(new_n1019), .B2(new_n821), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(new_n930), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1104), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1006), .B1(new_n1018), .B2(new_n1086), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1106), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1107), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT120), .B(new_n606), .C1(new_n1108), .C2(KEYINPUT60), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n930), .B(KEYINPUT120), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1104), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1107), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1996), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1042), .A2(new_n1048), .A3(new_n1002), .A4(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1018), .B2(new_n1006), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n549), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1132), .A3(new_n549), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(KEYINPUT59), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1099), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1129), .B2(new_n549), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT118), .B(new_n851), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1124), .A2(new_n1134), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1121), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n1124), .A4(new_n1136), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1116), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G2078), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1042), .A2(new_n1048), .A3(new_n1002), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1961), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1056), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1004), .A2(new_n486), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n634), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT123), .B(G2078), .Z(new_n1157));
  NOR4_X1   g732(.A1(new_n477), .A2(new_n1149), .A3(new_n1041), .A4(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1158), .A3(new_n1002), .A4(new_n1048), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1150), .A2(new_n1152), .A3(new_n1159), .ZN(new_n1160));
  OR3_X1    g735(.A1(new_n1160), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1149), .A2(new_n1148), .B1(new_n1056), .B2(new_n1151), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1149), .A2(G2078), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1075), .A2(new_n1076), .A3(new_n1048), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(G171), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n1160), .B2(G171), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1161), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1160), .A2(G171), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1162), .A2(G301), .A3(new_n1164), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT54), .ZN(new_n1173));
  AND4_X1   g748(.A1(new_n1093), .A2(new_n1173), .A3(new_n1069), .A4(new_n1039), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1048), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1002), .A2(G160), .A3(G40), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1073), .ZN(new_n1177));
  AOI21_X1  g752(.A(G1966), .B1(new_n1177), .B2(new_n1076), .ZN(new_n1178));
  OAI21_X1  g753(.A(G286), .B1(new_n1178), .B2(new_n1072), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1077), .A2(new_n749), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1072), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(G168), .A3(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1179), .A2(G8), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT121), .B1(new_n1078), .B2(new_n1020), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT51), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(G8), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(KEYINPUT51), .B2(new_n1184), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1170), .B(new_n1174), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1097), .B1(new_n1146), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1020), .B1(new_n1078), .B2(G168), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1179), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(KEYINPUT51), .A3(new_n1184), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1071), .A2(G171), .A3(new_n1093), .A4(new_n1165), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1016), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1007), .A2(new_n1125), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT46), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1007), .B1(new_n1008), .B2(new_n797), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT47), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n726), .A2(new_n728), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT125), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1010), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1208), .B1(new_n821), .B2(new_n819), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1012), .A2(KEYINPUT126), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1013), .A2(G1986), .A3(G290), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1213), .B1(new_n1012), .B2(KEYINPUT126), .ZN(new_n1214));
  OAI221_X1 g789(.A(new_n1205), .B1(new_n1209), .B2(new_n1013), .C1(new_n1210), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1200), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g792(.A(G401), .ZN(new_n1219));
  NOR2_X1   g793(.A1(G227), .A2(new_n459), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n1219), .A2(new_n696), .A3(new_n695), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g795(.A(new_n1221), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n994), .B(new_n1222), .C1(new_n912), .C2(new_n919), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


