//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143, new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT70), .Z(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n463), .B2(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT71), .B1(new_n469), .B2(new_n460), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n460), .B1(new_n473), .B2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n470), .B2(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n472), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n460), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n460), .C1(new_n471), .C2(new_n472), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT73), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(G138), .A3(new_n490), .A4(new_n460), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n506), .A2(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n513), .A2(new_n514), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n509), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n533), .A2(new_n510), .B1(new_n516), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n520), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n539), .A2(new_n510), .B1(new_n516), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n520), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT74), .Z(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  AND2_X1   g125(.A1(G78), .A2(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT77), .ZN(new_n552));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n513), .B2(new_n514), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(KEYINPUT76), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n509), .A2(G91), .A3(new_n515), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n558), .A2(new_n556), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n556), .B1(new_n558), .B2(KEYINPUT76), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  XNOR2_X1  g141(.A(G168), .B(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  NOR2_X1   g143(.A1(new_n507), .A2(new_n508), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n512), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n516), .ZN(G288));
  NAND2_X1  g149(.A1(new_n570), .A2(G48), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n575), .B1(new_n516), .B2(new_n576), .C1(new_n520), .C2(new_n577), .ZN(G305));
  NOR2_X1   g153(.A1(new_n528), .A2(new_n569), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G85), .B1(G47), .B2(new_n570), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT79), .Z(new_n581));
  AOI22_X1  g156(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n579), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  AOI22_X1  g162(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n520), .B1(new_n588), .B2(KEYINPUT80), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(KEYINPUT80), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n570), .A2(G54), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G321));
  XOR2_X1   g168(.A(G321), .B(KEYINPUT81), .Z(G284));
  NOR2_X1   g169(.A1(G299), .A2(G868), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n567), .B2(G868), .ZN(G297));
  AOI21_X1  g171(.A(new_n595), .B1(new_n567), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n592), .B1(new_n598), .B2(G860), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n598), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n463), .A2(new_n461), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n480), .A2(G135), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n482), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n460), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G2096), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n609), .A2(new_n610), .A3(new_n617), .ZN(G156));
  INV_X1    g193(.A(KEYINPUT14), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(G401));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT17), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2100), .Z(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(new_n616), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1971), .B(G1976), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1956), .B(G2474), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1961), .B(G1966), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT20), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n647), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n647), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1991), .B(G1996), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G229));
  INV_X1    g237(.A(G16), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G20), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT23), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(G299), .B2(G16), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1956), .ZN(new_n667));
  INV_X1    g242(.A(G29), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G33), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n480), .A2(G139), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n463), .A2(G127), .ZN(new_n677));
  AND2_X1   g252(.A1(G115), .A2(G2104), .ZN(new_n678));
  OAI21_X1  g253(.A(G2105), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n669), .B1(new_n680), .B2(new_n668), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G2072), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n504), .A2(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n668), .A2(G27), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G2084), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT24), .B(G34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(new_n668), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  INV_X1    g266(.A(G160), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n668), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n687), .A2(G2078), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G2078), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n681), .A2(G2072), .B1(new_n695), .B2(new_n686), .ZN(new_n696));
  AND4_X1   g271(.A1(new_n667), .A2(new_n683), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1961), .ZN(new_n698));
  NOR2_X1   g273(.A1(G171), .A2(new_n663), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G5), .B2(new_n663), .ZN(new_n700));
  NOR2_X1   g275(.A1(G168), .A2(new_n663), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n663), .B2(G21), .ZN(new_n702));
  INV_X1    g277(.A(G1966), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n698), .A2(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n668), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n461), .A2(G105), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n461), .A2(KEYINPUT95), .A3(G105), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n708), .A2(new_n709), .B1(new_n480), .B2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G129), .B2(new_n482), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n705), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G19), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n544), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT89), .B(G1341), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n704), .B1(new_n715), .B2(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n668), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT96), .B1(new_n615), .B2(new_n668), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n668), .B1(new_n724), .B2(G28), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT97), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(KEYINPUT97), .B1(new_n724), .B2(G28), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n700), .A2(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n720), .A2(new_n721), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n693), .A2(new_n688), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n718), .A2(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT29), .B(G2090), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n733), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n663), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n592), .B2(new_n663), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1348), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n668), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n482), .A2(G128), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n460), .A2(G116), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n749), .A2(KEYINPUT90), .A3(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(KEYINPUT90), .B1(new_n749), .B2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2067), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n742), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n697), .A2(new_n732), .A3(new_n739), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n663), .A2(G22), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G166), .B2(new_n663), .ZN(new_n757));
  INV_X1    g332(.A(G1971), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G23), .B(G288), .S(G16), .Z(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT33), .B(G1976), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT88), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G6), .A2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G48), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n765), .A2(new_n510), .B1(new_n516), .B2(new_n576), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n577), .A2(new_n520), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n764), .B1(new_n768), .B2(G16), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT32), .B(G1981), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n759), .A2(new_n763), .A3(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT34), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n663), .A2(G24), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT86), .Z(new_n775));
  INV_X1    g350(.A(G290), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n776), .A2(KEYINPUT87), .ZN(new_n777));
  OAI21_X1  g352(.A(G16), .B1(new_n776), .B2(KEYINPUT87), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G1986), .ZN(new_n780));
  NOR2_X1   g355(.A1(G25), .A2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G95), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n782), .A2(new_n460), .A3(KEYINPUT84), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT84), .B1(new_n782), .B2(new_n460), .ZN(new_n784));
  OAI221_X1 g359(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n480), .A2(G131), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n482), .A2(G119), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT85), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n790), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n779), .B2(G1986), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n773), .A2(new_n780), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT36), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT36), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n755), .B1(new_n796), .B2(new_n797), .ZN(G311));
  XNOR2_X1  g373(.A(G311), .B(KEYINPUT98), .ZN(G150));
  NAND2_X1  g374(.A1(new_n592), .A2(G559), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT38), .ZN(new_n801));
  NAND2_X1  g376(.A1(G80), .A2(G543), .ZN(new_n802));
  INV_X1    g377(.A(G67), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n528), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n520), .B1(new_n804), .B2(KEYINPUT99), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT99), .B2(new_n804), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n579), .A2(G93), .B1(G55), .B2(new_n570), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n544), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n806), .A2(new_n544), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n801), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT100), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n808), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  INV_X1    g395(.A(G37), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n714), .B(new_n749), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n680), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n500), .B1(new_n493), .B2(new_n492), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n482), .A2(G130), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n460), .A2(G118), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G142), .B2(new_n480), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(new_n606), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n788), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n825), .A2(new_n832), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n615), .B(new_n486), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n692), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n833), .A2(new_n834), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n836), .A2(new_n833), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n821), .B1(new_n840), .B2(new_n841), .C1(new_n839), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g419(.A(G290), .B(G305), .ZN(new_n845));
  XNOR2_X1  g420(.A(G303), .B(G288), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G290), .B(new_n768), .ZN(new_n848));
  INV_X1    g423(.A(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT42), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n847), .A2(new_n850), .A3(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n851), .B1(new_n856), .B2(KEYINPUT42), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n592), .A2(G299), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n564), .A3(new_n561), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(KEYINPUT102), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n592), .A2(new_n862), .A3(G299), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(KEYINPUT41), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n858), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n863), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n601), .B(new_n812), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n867), .B(new_n868), .S(new_n869), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n857), .B(new_n870), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n808), .B(new_n871), .S(G868), .Z(G295));
  MUX2_X1   g447(.A(new_n808), .B(new_n871), .S(G868), .Z(G331));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n874));
  NOR2_X1   g449(.A1(G171), .A2(G168), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n567), .B2(G171), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(new_n812), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n812), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n863), .A3(new_n861), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n864), .A2(new_n866), .A3(new_n877), .A4(new_n878), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n854), .A2(new_n855), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n821), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n854), .A2(new_n855), .B1(new_n881), .B2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n874), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n868), .B1(new_n879), .B2(new_n865), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n858), .A2(new_n860), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT41), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n855), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT103), .B1(new_n850), .B2(new_n847), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n886), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n821), .A3(new_n882), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n885), .B1(new_n874), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT44), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n891), .A2(new_n882), .A3(new_n874), .A4(new_n821), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n883), .B2(new_n884), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n895), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n899), .B2(KEYINPUT104), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n894), .B1(new_n900), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g476(.A(new_n500), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n494), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G1384), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n480), .A2(G137), .B1(G101), .B2(new_n461), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n474), .A2(new_n475), .ZN(new_n909));
  AOI211_X1 g484(.A(KEYINPUT71), .B(new_n460), .C1(new_n473), .C2(new_n467), .ZN(new_n910));
  OAI211_X1 g485(.A(G40), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT106), .Z(new_n913));
  INV_X1    g488(.A(G1996), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n915), .A2(KEYINPUT46), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(KEYINPUT46), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n749), .B(G2067), .Z(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n713), .A3(new_n710), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n916), .A2(new_n917), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n714), .B(new_n914), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n789), .A2(new_n791), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n789), .A2(new_n791), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n913), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1986), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n913), .A2(new_n928), .A3(new_n776), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT126), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n931), .B2(KEYINPUT48), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(KEYINPUT48), .B2(new_n931), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n923), .A2(new_n925), .B1(G2067), .B2(new_n749), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n921), .B(new_n933), .C1(new_n913), .C2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n906), .A2(G1384), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n504), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT109), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n504), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(G40), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n941), .B(new_n466), .C1(new_n470), .C2(new_n476), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n905), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n940), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n504), .B2(new_n904), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n824), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(new_n911), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n945), .A2(new_n703), .B1(new_n949), .B2(new_n688), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT51), .B1(new_n950), .B2(G168), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n911), .ZN(new_n952));
  INV_X1    g527(.A(new_n947), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n688), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n494), .B2(new_n902), .ZN(new_n955));
  OAI211_X1 g530(.A(G160), .B(G40), .C1(KEYINPUT45), .C2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n504), .A2(new_n939), .A3(new_n936), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n939), .B1(new_n504), .B2(new_n936), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(G168), .B(new_n954), .C1(new_n959), .C2(G1966), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G8), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n960), .B2(G8), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT119), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n966), .B(new_n967), .C1(new_n961), .C2(new_n951), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT124), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n964), .A2(new_n968), .A3(new_n971), .A4(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n952), .A2(new_n953), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n698), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n959), .A2(KEYINPUT53), .A3(new_n695), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n943), .B(G1384), .C1(new_n494), .C2(new_n902), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(new_n911), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n504), .A2(new_n904), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n906), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n695), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT121), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n975), .B(new_n976), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G171), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT122), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT122), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n989), .A3(G171), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G303), .A2(G8), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT55), .Z(new_n993));
  INV_X1    g568(.A(new_n906), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n504), .B2(new_n904), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n995), .A2(new_n911), .A3(new_n977), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G1971), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n974), .A2(G2090), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n993), .B(G8), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n911), .A2(new_n905), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1001), .B(new_n1002), .C1(new_n1004), .C2(KEYINPUT49), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  OAI221_X1 g587(.A(G8), .B1(new_n1012), .B2(G288), .C1(new_n911), .C2(new_n905), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1012), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1011), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n999), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n504), .A2(new_n946), .A3(new_n904), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT50), .B1(new_n824), .B2(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n942), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n996), .A2(G1971), .B1(new_n1022), .B2(G2090), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n993), .B1(G8), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n991), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT62), .B1(new_n964), .B2(new_n968), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT125), .B1(new_n973), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n949), .A2(G1348), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n911), .A2(new_n905), .A3(G2067), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n592), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT56), .B(G2072), .ZN(new_n1035));
  INV_X1    g610(.A(G1956), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n996), .A2(new_n1035), .B1(new_n1022), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n561), .A2(new_n1038), .A3(new_n1039), .A4(new_n564), .ZN(new_n1040));
  NAND2_X1  g615(.A1(KEYINPUT111), .A2(KEYINPUT57), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  INV_X1    g617(.A(new_n564), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1041), .B(new_n1042), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1022), .A2(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n978), .A2(new_n980), .A3(new_n1035), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1048), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1034), .A2(new_n1047), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT112), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n978), .A2(new_n980), .A3(new_n1035), .ZN(new_n1057));
  AND4_X1   g632(.A1(KEYINPUT112), .A2(new_n1046), .A3(new_n1050), .A4(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1047), .A2(new_n1064), .A3(new_n1053), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT118), .ZN(new_n1066));
  NOR4_X1   g641(.A1(new_n1031), .A2(KEYINPUT60), .A3(new_n859), .A4(new_n1032), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1032), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n859), .C1(new_n949), .C2(G1348), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1033), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(KEYINPUT60), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1047), .A2(new_n1064), .A3(new_n1053), .A4(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1063), .A2(new_n1066), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NOR4_X1   g650(.A1(new_n995), .A2(new_n977), .A3(new_n911), .A4(G1996), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n911), .B2(new_n905), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n978), .A2(new_n914), .A3(new_n980), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1078), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n809), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1081), .A2(new_n1082), .A3(new_n1078), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1082), .B1(new_n1081), .B2(new_n1078), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n544), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1085), .B(new_n544), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT117), .A3(new_n1085), .A4(new_n544), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1086), .A2(new_n1090), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1059), .B1(new_n1074), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT123), .B(G2078), .Z(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n466), .A2(new_n474), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n907), .B(new_n1101), .C1(new_n943), .C2(new_n905), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n975), .B(new_n1102), .C1(new_n984), .C2(new_n985), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1098), .B1(new_n991), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(G171), .ZN(new_n1106));
  NOR4_X1   g681(.A1(new_n995), .A2(new_n977), .A3(new_n911), .A4(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(new_n983), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(G301), .A3(new_n975), .A4(new_n976), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(KEYINPUT54), .A3(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n964), .A2(new_n1113), .A3(new_n968), .A4(new_n1025), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1097), .A2(new_n1105), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1018), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1009), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G288), .A2(G1976), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1011), .A2(new_n1118), .B1(new_n1000), .B2(new_n768), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1116), .A2(new_n999), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n950), .A2(new_n1008), .A3(G286), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT110), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1019), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n998), .B2(new_n997), .ZN(new_n1126));
  INV_X1    g701(.A(new_n993), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1125), .B1(new_n1130), .B2(new_n1122), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1120), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1029), .A2(new_n1030), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n929), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n776), .A2(new_n928), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n913), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT107), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n927), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n935), .B1(new_n1134), .B2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g715(.A(G227), .ZN(new_n1142));
  NAND2_X1  g716(.A1(G319), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g717(.A1(G229), .A2(G401), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g718(.A1(new_n843), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g719(.A1(new_n900), .A2(new_n1145), .ZN(G308));
  OR2_X1    g720(.A1(new_n900), .A2(new_n1145), .ZN(G225));
endmodule


