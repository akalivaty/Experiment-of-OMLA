//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n206), .B1(G155gat), .B2(G162gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n208), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n208), .A2(new_n218), .A3(KEYINPUT74), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G127gat), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G113gat), .ZN(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n208), .A2(new_n218), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n208), .A2(new_n218), .A3(KEYINPUT75), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n239), .A3(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n250), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT4), .B1(new_n241), .B2(new_n240), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n256), .A2(KEYINPUT77), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT77), .B1(new_n256), .B2(new_n257), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n243), .B(new_n246), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n241), .B(new_n240), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n245), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n241), .A2(new_n240), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n243), .B2(KEYINPUT4), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT75), .B1(new_n208), .B2(new_n218), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n208), .A2(new_n218), .A3(KEYINPUT75), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n231), .A2(new_n239), .A3(KEYINPUT67), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n231), .B2(new_n239), .ZN(new_n268));
  OAI22_X1  g067(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n244), .B1(new_n269), .B2(new_n255), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT5), .B(new_n262), .C1(new_n264), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n260), .B2(new_n271), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n278), .B(new_n276), .C1(new_n260), .C2(new_n271), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  AND3_X1   g083(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n286), .A2(new_n287), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(new_n290), .A3(new_n297), .A4(new_n291), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n301), .A2(G169gat), .A3(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(G169gat), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n302), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n299), .A3(new_n300), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n311), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n295), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n290), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT25), .ZN(new_n316));
  AND2_X1   g115(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n295), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT26), .ZN(new_n321));
  OR3_X1    g120(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n306), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n295), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n320), .A2(new_n323), .A3(new_n326), .A4(new_n288), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n316), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n316), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT29), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n300), .B1(new_n308), .B2(new_n314), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n320), .A2(new_n326), .A3(new_n288), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n323), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n333), .A3(new_n309), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT22), .ZN(new_n342));
  INV_X1    g141(.A(G211gat), .ZN(new_n343));
  INV_X1    g142(.A(G218gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G211gat), .B(G218gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT68), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n341), .A3(new_n345), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(KEYINPUT68), .A3(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n330), .B1(new_n338), .B2(new_n309), .ZN(new_n357));
  INV_X1    g156(.A(new_n331), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n333), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n354), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n328), .A2(new_n334), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G8gat), .B(G36gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(G92gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT71), .B(G64gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  NAND3_X1  g167(.A1(new_n356), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n364), .A3(KEYINPUT72), .A4(new_n368), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n356), .A2(new_n364), .A3(KEYINPUT30), .A4(new_n368), .ZN(new_n375));
  INV_X1    g174(.A(new_n368), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n332), .B1(new_n329), .B2(new_n331), .ZN(new_n377));
  INV_X1    g176(.A(new_n363), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n377), .A2(new_n361), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n354), .B1(new_n335), .B2(new_n339), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n283), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT79), .B(G22gat), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n241), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g187(.A(G228gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n222), .B2(new_n223), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n388), .B(new_n391), .C1(new_n361), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n349), .B2(new_n351), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n219), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n250), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n392), .A2(new_n355), .ZN(new_n400));
  OAI22_X1  g199(.A1(new_n399), .A2(new_n400), .B1(new_n389), .B2(new_n390), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n386), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n401), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT80), .B1(new_n409), .B2(new_n385), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n404), .B(new_n408), .C1(new_n410), .C2(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(G22gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n407), .C1(new_n409), .C2(new_n385), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n338), .A2(new_n254), .A3(new_n309), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n267), .A2(new_n268), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n328), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G227gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n390), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT32), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n420), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n415), .B2(new_n417), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT32), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT34), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n418), .A2(new_n420), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n423), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n423), .B2(new_n427), .ZN(new_n431));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n425), .B2(KEYINPUT33), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n430), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n422), .B1(new_n421), .B2(KEYINPUT32), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT34), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n428), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n427), .A3(new_n429), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n384), .A2(KEYINPUT35), .A3(new_n414), .A4(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n374), .A2(new_n382), .ZN(new_n445));
  INV_X1    g244(.A(new_n280), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n278), .A3(new_n277), .ZN(new_n447));
  INV_X1    g246(.A(new_n282), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n445), .A2(new_n443), .A3(new_n449), .A4(new_n414), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(new_n449), .ZN(new_n454));
  INV_X1    g253(.A(new_n414), .ZN(new_n455));
  INV_X1    g254(.A(new_n442), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n437), .A3(new_n441), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT36), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n436), .B2(new_n442), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n454), .A2(new_n455), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n261), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT81), .B1(new_n261), .B2(new_n245), .ZN(new_n465));
  INV_X1    g264(.A(new_n243), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n257), .B1(new_n269), .B2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n256), .A2(KEYINPUT77), .A3(new_n257), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n464), .B(new_n465), .C1(new_n471), .C2(new_n244), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n243), .B1(new_n258), .B2(new_n259), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n463), .A3(new_n245), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(KEYINPUT40), .A3(new_n276), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n276), .A3(new_n474), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n383), .A2(new_n446), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n356), .A2(new_n364), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n376), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT38), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n361), .B1(new_n377), .B2(new_n378), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT83), .B(new_n361), .C1(new_n377), .C2(new_n378), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n489), .B(new_n490), .C1(new_n355), .C2(new_n340), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT37), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n371), .A2(new_n373), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT38), .B1(new_n495), .B2(new_n485), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n283), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n374), .A2(new_n382), .B1(new_n476), .B2(new_n477), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n475), .A2(new_n446), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n481), .A2(new_n414), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n453), .B1(new_n461), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G230gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n390), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n506));
  INV_X1    g305(.A(G85gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(G85gat), .A3(G92gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n509), .A2(new_n511), .B1(KEYINPUT8), .B2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G99gat), .B(G106gat), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT93), .B(G92gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n513), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n506), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n513), .A2(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT95), .A3(new_n518), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n524), .B(new_n525), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n531), .B(new_n506), .C1(new_n519), .C2(new_n520), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT10), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n519), .B2(new_n520), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(KEYINPUT94), .A3(new_n518), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n536), .A4(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n505), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n530), .A2(new_n504), .A3(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G120gat), .B(G148gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n546));
  INV_X1    g345(.A(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n539), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n536), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(KEYINPUT86), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT86), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G29gat), .A2(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n563), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n567), .B2(new_n559), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT15), .A3(new_n556), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n553), .B(new_n555), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  AND4_X1   g369(.A1(KEYINPUT86), .A2(new_n566), .A3(new_n552), .A4(new_n569), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n551), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n569), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n535), .A2(new_n573), .A3(new_n536), .ZN(new_n574));
  NAND3_X1  g373(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT92), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n577), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n572), .A2(new_n583), .A3(new_n574), .A4(new_n575), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n578), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n502), .A2(new_n550), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G211gat), .ZN(new_n590));
  INV_X1    g389(.A(G15gat), .ZN(new_n591));
  INV_X1    g390(.A(G22gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G15gat), .A2(G22gat), .ZN(new_n594));
  INV_X1    g393(.A(G1gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n593), .A2(new_n594), .B1(KEYINPUT16), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n594), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(G1gat), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(G8gat), .B1(new_n600), .B2(KEYINPUT88), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT87), .A3(G8gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n599), .A2(G1gat), .ZN(new_n603));
  OAI21_X1  g402(.A(G8gat), .B1(new_n603), .B2(new_n596), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n597), .A2(new_n601), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G183gat), .ZN(new_n610));
  INV_X1    g409(.A(G231gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n390), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n609), .B(new_n294), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n612), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n590), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT91), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n610), .A2(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n612), .ZN(new_n623));
  INV_X1    g422(.A(new_n590), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n617), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n621), .B1(new_n617), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n607), .B1(new_n570), .B2(new_n571), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT88), .B1(new_n603), .B2(new_n596), .ZN(new_n632));
  INV_X1    g431(.A(G8gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n597), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT87), .B1(new_n600), .B2(G8gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n604), .A2(new_n605), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n573), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G113gat), .B(G141gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G197gat), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT11), .B(G169gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  INV_X1    g445(.A(new_n573), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n607), .A2(KEYINPUT89), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT89), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n637), .B2(new_n573), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n650), .A3(new_n638), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n631), .B(KEYINPUT13), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n630), .A2(KEYINPUT18), .A3(new_n631), .A4(new_n638), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n641), .A2(new_n646), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n653), .A3(new_n654), .ZN(new_n658));
  INV_X1    g457(.A(new_n646), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n629), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n588), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n449), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n595), .ZN(G1324gat));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n445), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  OR2_X1    g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT42), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n671), .A2(new_n633), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n458), .A2(new_n460), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n668), .A2(new_n591), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n588), .A2(new_n667), .A3(new_n443), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n591), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n668), .A2(new_n414), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n592), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT98), .B(KEYINPUT43), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n587), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n501), .A2(new_n461), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n450), .B(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n666), .A2(new_n628), .A3(new_n550), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n449), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n690), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n691), .B(KEYINPUT99), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n449), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(G1328gat));
  OR3_X1    g499(.A1(new_n698), .A2(KEYINPUT100), .A3(new_n445), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT100), .B1(new_n698), .B2(new_n445), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(G36gat), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n692), .A2(G36gat), .A3(new_n445), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(new_n443), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n692), .A2(G43gat), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n679), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n696), .A2(new_n709), .A3(new_n697), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n710), .B2(G43gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g511(.A1(new_n455), .A2(G50gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n692), .A2(new_n414), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n698), .A2(new_n713), .B1(G50gat), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g515(.A(new_n550), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n657), .A2(new_n660), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n662), .A2(new_n663), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n587), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n628), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n502), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n283), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT101), .B(G57gat), .Z(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  NAND2_X1  g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n383), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT102), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  INV_X1    g529(.A(new_n722), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n731), .A2(G71gat), .A3(new_n707), .ZN(new_n732));
  OAI21_X1  g531(.A(G71gat), .B1(new_n731), .B2(new_n679), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n455), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n628), .A2(new_n665), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n502), .A2(KEYINPUT51), .A3(new_n687), .A4(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n690), .B2(new_n738), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(new_n742), .A3(new_n717), .ZN(new_n743));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743), .B2(new_n283), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n550), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT103), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n696), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n449), .A2(new_n507), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(new_n516), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(new_n383), .A3(new_n752), .A4(new_n746), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n679), .B1(new_n384), .B2(new_n414), .ZN(new_n759));
  INV_X1    g558(.A(new_n500), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT82), .B1(new_n498), .B2(new_n499), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n497), .A2(new_n414), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n587), .B(new_n738), .C1(new_n764), .C2(new_n453), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n690), .A2(new_n741), .A3(new_n738), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n445), .A2(G92gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n550), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n757), .A2(new_n758), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n740), .A2(new_n742), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(KEYINPUT104), .A3(new_n550), .A4(new_n768), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n750), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n778), .A2(KEYINPUT105), .A3(KEYINPUT52), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT105), .B1(new_n778), .B2(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n743), .A2(new_n782), .A3(new_n443), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n747), .A2(new_n709), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(G1338gat));
  NAND2_X1  g584(.A1(new_n743), .A2(new_n455), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n747), .A2(G106gat), .A3(new_n455), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT53), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n628), .A2(new_n720), .A3(new_n717), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n651), .A2(new_n652), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n631), .B1(new_n630), .B2(new_n638), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n645), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n655), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n655), .B2(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n587), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n530), .A2(new_n532), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n504), .B(new_n537), .C1(new_n805), .C2(KEYINPUT10), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(new_n539), .A3(KEYINPUT54), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n505), .C1(new_n533), .C2(new_n538), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n544), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n539), .A3(KEYINPUT54), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n544), .A4(new_n809), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(new_n549), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n803), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n655), .A2(new_n799), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n550), .B1(new_n585), .B2(new_n586), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n815), .A2(new_n720), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n796), .B1(new_n629), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n795), .B1(new_n819), .B2(new_n455), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n449), .A2(new_n383), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n628), .A2(new_n720), .A3(new_n717), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n817), .A2(new_n816), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n549), .A3(new_n813), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n655), .A2(new_n799), .A3(new_n800), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n587), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n687), .B1(new_n661), .B2(new_n664), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n822), .B1(new_n830), .B2(new_n628), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(KEYINPUT109), .A3(new_n414), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n820), .A2(new_n443), .A3(new_n821), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n666), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n455), .A3(new_n707), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n821), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n665), .A2(new_n234), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT110), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n833), .B2(new_n717), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n550), .A2(new_n232), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT111), .Z(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n836), .B2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n833), .A2(new_n227), .A3(new_n629), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n836), .A2(KEYINPUT112), .A3(new_n629), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT112), .B1(new_n836), .B2(new_n629), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n227), .ZN(G1342gat));
  OR3_X1    g647(.A1(new_n687), .A2(new_n383), .A3(KEYINPUT113), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT113), .B1(new_n687), .B2(new_n383), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n283), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n225), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n833), .B2(new_n687), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT114), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n455), .ZN(new_n859));
  INV_X1    g658(.A(new_n821), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n709), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n665), .A2(new_n211), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(KEYINPUT117), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  INV_X1    g669(.A(new_n868), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n830), .B2(new_n628), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n818), .A2(new_n629), .A3(KEYINPUT115), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n822), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n414), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n878), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n709), .A2(new_n860), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n665), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n882), .A2(KEYINPUT118), .A3(new_n665), .A4(new_n883), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(G141gat), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT58), .B1(new_n867), .B2(new_n868), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n861), .A2(new_n209), .A3(new_n550), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n883), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n717), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n209), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n831), .A2(KEYINPUT57), .A3(new_n455), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n859), .A2(new_n903), .A3(new_n878), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n902), .A2(new_n550), .A3(new_n883), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n897), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n900), .B2(new_n906), .ZN(G1345gat));
  NOR3_X1   g706(.A1(new_n898), .A2(new_n215), .A3(new_n629), .ZN(new_n908));
  AOI21_X1  g707(.A(G155gat), .B1(new_n861), .B2(new_n628), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n898), .B2(new_n687), .ZN(new_n911));
  OR4_X1    g710(.A1(G162gat), .A2(new_n859), .A3(new_n709), .A4(new_n851), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n445), .A2(new_n283), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n835), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n303), .A3(new_n665), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n820), .A2(new_n443), .A3(new_n832), .A4(new_n914), .ZN(new_n918));
  OAI21_X1  g717(.A(G169gat), .B1(new_n918), .B2(new_n666), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n304), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n550), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT121), .B1(new_n921), .B2(new_n550), .ZN(new_n923));
  AOI21_X1  g722(.A(G176gat), .B1(new_n916), .B2(new_n550), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(G1349gat));
  NAND3_X1  g724(.A1(new_n916), .A2(new_n628), .A3(new_n324), .ZN(new_n926));
  OAI21_X1  g725(.A(G183gat), .B1(new_n918), .B2(new_n629), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1350gat));
  NOR3_X1   g729(.A1(new_n915), .A2(G190gat), .A3(new_n687), .ZN(new_n931));
  OAI21_X1  g730(.A(G190gat), .B1(new_n918), .B2(new_n687), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(G190gat), .C1(new_n918), .C2(new_n687), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1351gat));
  XNOR2_X1  g737(.A(KEYINPUT124), .B(G197gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n914), .A2(new_n679), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n902), .A2(new_n904), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n942), .B2(new_n666), .ZN(new_n943));
  INV_X1    g742(.A(new_n940), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n831), .A2(new_n455), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n666), .B2(new_n946), .ZN(G1352gat));
  OR2_X1    g746(.A1(new_n945), .A2(G204gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n948), .A2(new_n717), .B1(new_n949), .B2(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND4_X1  g751(.A1(new_n902), .A2(new_n550), .A3(new_n904), .A4(new_n941), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  OR3_X1    g754(.A1(new_n945), .A2(G211gat), .A3(new_n629), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n902), .A2(new_n628), .A3(new_n904), .A4(new_n944), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g761(.A(KEYINPUT127), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1354gat));
  NOR3_X1   g763(.A1(new_n942), .A2(new_n344), .A3(new_n687), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n945), .A2(new_n687), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n344), .B2(new_n966), .ZN(G1355gat));
endmodule


