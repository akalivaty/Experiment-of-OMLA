//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(KEYINPUT11), .C1(new_n197), .C2(G137), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT11), .B1(new_n203), .B2(new_n199), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n201), .B2(new_n204), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n196), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT66), .B1(new_n214), .B2(G116), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n212), .A3(G119), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n219), .A2(new_n220), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n218), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n190), .A3(new_n192), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n191), .A2(KEYINPUT1), .A3(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n225), .B(new_n226), .C1(G128), .C2(new_n194), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n203), .A2(new_n198), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n210), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n211), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n196), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n199), .B1(new_n197), .B2(G137), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n200), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n207), .B1(new_n237), .B2(new_n198), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n208), .B1(new_n236), .B2(new_n200), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n233), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n222), .A4(new_n230), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G101), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n243), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n232), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n232), .A2(KEYINPUT69), .A3(new_n242), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n214), .A2(G116), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n216), .B1(new_n212), .B2(G119), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n214), .A2(KEYINPUT66), .A3(G116), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n221), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT2), .A2(G113), .ZN(new_n260));
  INV_X1    g074(.A(new_n220), .ZN(new_n261));
  NAND3_X1  g075(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n218), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n239), .B1(new_n205), .B2(G131), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n266), .B(new_n230), .C1(new_n267), .C2(new_n196), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n240), .B2(new_n230), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n254), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n188), .B1(new_n253), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n251), .A2(new_n252), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n271), .A4(new_n254), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n230), .B1(new_n267), .B2(new_n196), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n265), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n232), .A2(new_n278), .A3(new_n242), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n240), .A2(new_n222), .A3(new_n230), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n250), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n276), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n288), .B(new_n285), .C1(new_n273), .C2(new_n275), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT71), .B(new_n187), .C1(new_n287), .C2(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n187), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n273), .A2(new_n275), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n288), .B1(new_n297), .B2(new_n285), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n276), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n283), .B1(new_n279), .B2(KEYINPUT28), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT29), .A3(new_n250), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n249), .B(new_n283), .C1(new_n279), .C2(KEYINPUT28), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT72), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n301), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n271), .A2(new_n232), .A3(new_n242), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n249), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  INV_X1    g127(.A(new_n303), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n249), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n307), .A2(KEYINPUT72), .A3(KEYINPUT29), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n305), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT73), .A4(new_n302), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n309), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n300), .A2(KEYINPUT32), .B1(new_n319), .B2(G472), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n295), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G234), .ZN(new_n322));
  OAI21_X1  g136(.A(G217), .B1(new_n322), .B2(G902), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT74), .Z(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G119), .B(G128), .Z(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n214), .B2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n330), .B(new_n331), .C1(G119), .C2(new_n223), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(G110), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G125), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT75), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n334), .A2(KEYINPUT75), .A3(G125), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n340), .A2(new_n189), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n189), .B1(new_n340), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n333), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n333), .B(new_n347), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n326), .A2(new_n327), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n332), .B2(G110), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n335), .A2(new_n337), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n189), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(new_n344), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n245), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT77), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n349), .A2(new_n356), .A3(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(new_n365), .B2(new_n302), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n361), .B1(new_n349), .B2(new_n356), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n355), .B(new_n362), .C1(new_n346), .C2(new_n348), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n302), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n325), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n323), .A2(new_n302), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n302), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n370), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n324), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT78), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n267), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT79), .B(G101), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT3), .A3(G104), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT3), .B1(new_n389), .B2(G104), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n386), .B(new_n388), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n389), .B2(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(G104), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(KEYINPUT80), .A3(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n226), .B1(new_n194), .B2(G128), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n401), .A2(new_n402), .B1(new_n194), .B2(new_n224), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT81), .B(new_n226), .C1(new_n194), .C2(G128), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n387), .B2(G107), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(new_n390), .B1(new_n387), .B2(G107), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n408), .A2(new_n386), .B1(new_n398), .B2(G101), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n227), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT12), .B(new_n385), .C1(new_n405), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n385), .B1(new_n405), .B2(new_n410), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G128), .B1(new_n190), .B2(new_n192), .ZN(new_n417));
  INV_X1    g231(.A(new_n226), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n225), .A3(new_n404), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n409), .ZN(new_n421));
  INV_X1    g235(.A(new_n401), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n400), .A2(new_n422), .A3(new_n225), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n267), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT82), .A3(KEYINPUT12), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT10), .B1(new_n420), .B2(new_n409), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n409), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n429));
  INV_X1    g243(.A(G101), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n408), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n196), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n393), .B(KEYINPUT4), .C1(new_n430), .C2(new_n408), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(new_n267), .A3(new_n429), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  INV_X1    g252(.A(G227), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G953), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n431), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n432), .A3(G101), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n233), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n429), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n427), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n448), .B2(new_n267), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n385), .B1(new_n447), .B2(new_n427), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n437), .A2(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G469), .B1(new_n451), .B2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n426), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n436), .A2(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n441), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT83), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n426), .A2(new_n449), .B1(new_n454), .B2(new_n441), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n460));
  NOR4_X1   g274(.A1(new_n459), .A2(new_n460), .A3(G469), .A4(G902), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n452), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT9), .B(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT84), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT5), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G113), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n409), .A3(new_n264), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT87), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n409), .A3(new_n473), .A4(new_n264), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n264), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n400), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT8), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n434), .A2(new_n265), .A3(new_n445), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n434), .A2(new_n265), .A3(new_n483), .A4(new_n445), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(new_n478), .A3(new_n471), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n227), .A2(new_n336), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n336), .B2(new_n196), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n245), .A2(G224), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(new_n302), .ZN(new_n492));
  INV_X1    g306(.A(new_n478), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n471), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n264), .A2(new_n259), .B1(new_n431), .B2(new_n432), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n483), .B1(new_n495), .B2(new_n434), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n488), .B(KEYINPUT86), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n487), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(new_n493), .C1(new_n494), .C2(new_n496), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n492), .B(new_n503), .C1(KEYINPUT88), .C2(new_n506), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n467), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n244), .A2(new_n245), .A3(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n191), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n244), .A2(new_n245), .A3(G143), .A4(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT17), .A3(G131), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n343), .A2(new_n344), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n516), .B(G131), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n519), .B(new_n520), .C1(KEYINPUT17), .C2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n387), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n514), .B(new_n515), .C1(new_n525), .C2(new_n207), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT90), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n516), .A2(KEYINPUT18), .A3(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n338), .A2(new_n339), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n353), .B(KEYINPUT89), .C1(new_n529), .C2(new_n189), .ZN(new_n530));
  OR3_X1    g344(.A1(new_n529), .A2(KEYINPUT89), .A3(new_n189), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n522), .A2(new_n524), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n344), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n352), .A2(KEYINPUT19), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n529), .B2(KEYINPUT19), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n521), .B(new_n534), .C1(G146), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n524), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G475), .A2(G902), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT92), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n512), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n512), .A3(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n223), .A2(G143), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n191), .A2(G128), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n197), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n212), .A2(KEYINPUT14), .A3(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(G116), .B(G122), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(G107), .B(new_n552), .C1(new_n554), .C2(KEYINPUT14), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n551), .B(new_n555), .C1(G107), .C2(new_n554), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n548), .A2(KEYINPUT13), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(new_n549), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n548), .A2(KEYINPUT13), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n197), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n553), .B(new_n389), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n550), .A2(new_n197), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n556), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G217), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n463), .A2(new_n565), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n556), .B(new_n566), .C1(new_n560), .C2(new_n563), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n302), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n573), .B(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n245), .A2(G952), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n322), .B2(new_n244), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n302), .B(new_n245), .C1(G234), .C2(G237), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT21), .B(G898), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n533), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n524), .B1(new_n522), .B2(new_n532), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n302), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G475), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n547), .A2(new_n577), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n465), .A2(new_n511), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n321), .A2(new_n384), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n386), .B(KEYINPUT94), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G3));
  AND4_X1   g407(.A1(new_n382), .A2(new_n377), .A3(new_n462), .A4(new_n464), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n302), .B1(new_n287), .B2(new_n289), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n594), .A2(new_n292), .A3(new_n294), .A4(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n546), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n588), .B1(new_n599), .B2(new_n544), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n573), .A2(new_n574), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n571), .A2(new_n572), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n568), .A2(KEYINPUT33), .A3(new_n570), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n302), .A2(G478), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(new_n584), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n467), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n504), .A2(new_n507), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n506), .B1(new_n492), .B2(new_n503), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n600), .ZN(new_n618));
  INV_X1    g432(.A(new_n577), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n584), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n613), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  AND2_X1   g439(.A1(new_n292), .A2(new_n294), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n462), .A2(new_n510), .A3(new_n464), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n357), .B(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n629), .A2(new_n375), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n380), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n589), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n626), .A2(new_n627), .A3(new_n596), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(new_n465), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n618), .A2(new_n619), .ZN(new_n637));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n581), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n579), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n613), .A2(new_n631), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n321), .A2(new_n636), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  NAND2_X1  g459(.A1(new_n508), .A2(new_n509), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT38), .Z(new_n647));
  INV_X1    g461(.A(new_n631), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n619), .A2(new_n600), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n647), .A2(new_n467), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n640), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n274), .A2(new_n271), .A3(new_n254), .ZN(new_n655));
  INV_X1    g469(.A(new_n279), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n250), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n657), .B2(new_n302), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n300), .B2(KEYINPUT32), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n295), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n650), .A2(new_n653), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n600), .A2(new_n608), .A3(new_n640), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n465), .A2(new_n613), .A3(new_n631), .A4(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n321), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n664), .B1(new_n321), .B2(new_n666), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  NAND2_X1  g484(.A1(new_n453), .A2(new_n455), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n457), .A3(new_n302), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n460), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n456), .A2(KEYINPUT83), .A3(new_n457), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n459), .B2(G902), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n464), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n321), .A2(new_n384), .A3(new_n614), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n321), .A2(new_n384), .A3(new_n621), .A4(new_n678), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  INV_X1    g497(.A(new_n613), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n678), .A2(new_n684), .A3(new_n632), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n295), .B2(new_n320), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n214), .ZN(G21));
  NAND2_X1  g501(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n595), .A2(new_n689), .A3(G472), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n380), .A2(new_n381), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n249), .B1(new_n303), .B2(KEYINPUT98), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(KEYINPUT98), .B2(new_n303), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n187), .B1(new_n694), .B2(new_n297), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n677), .A2(new_n583), .A3(new_n613), .A4(new_n649), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n692), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT100), .B(G122), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G24));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n595), .A2(new_n689), .A3(G472), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n689), .B1(new_n595), .B2(G472), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n648), .B(new_n695), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n677), .A2(new_n613), .ZN(new_n704));
  INV_X1    g518(.A(new_n665), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n700), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n695), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n688), .B2(new_n690), .ZN(new_n709));
  INV_X1    g523(.A(new_n706), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT101), .A4(new_n648), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NAND2_X1  g527(.A1(new_n462), .A2(KEYINPUT102), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n452), .B(new_n715), .C1(new_n458), .C2(new_n461), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n464), .A2(new_n508), .A3(new_n610), .A4(new_n509), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n714), .A2(new_n705), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n309), .A2(new_n315), .A3(new_n318), .ZN(new_n721));
  OAI22_X1  g535(.A1(new_n721), .A2(new_n654), .B1(new_n290), .B2(new_n293), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n290), .A2(new_n293), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n692), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n320), .A2(new_n723), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n692), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n720), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n383), .B1(new_n295), .B2(new_n320), .ZN(new_n731));
  INV_X1    g545(.A(new_n718), .ZN(new_n732));
  AOI211_X1 g546(.A(KEYINPUT103), .B(KEYINPUT42), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n321), .A2(new_n384), .A3(new_n732), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n719), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n730), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(KEYINPUT105), .B(new_n730), .C1(new_n733), .C2(new_n736), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n207), .ZN(G33));
  AND4_X1   g556(.A1(new_n642), .A2(new_n714), .A3(new_n716), .A4(new_n717), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n731), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT106), .B(G134), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G36));
  AOI21_X1  g560(.A(new_n631), .B1(new_n626), .B2(new_n596), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT109), .Z(new_n748));
  NAND2_X1  g562(.A1(new_n618), .A2(new_n608), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(KEYINPUT43), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT108), .Z(new_n755));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n646), .A2(new_n467), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n451), .A2(KEYINPUT45), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n451), .B2(KEYINPUT45), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n675), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n464), .A3(new_n651), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n756), .A2(new_n758), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n748), .A2(KEYINPUT44), .A3(new_n755), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT110), .B(G137), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G39));
  NAND2_X1  g586(.A1(new_n766), .A2(new_n464), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT47), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n383), .A2(new_n705), .A3(new_n757), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n774), .A2(new_n321), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n334), .ZN(G42));
  NAND2_X1  g591(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n728), .A2(new_n727), .A3(new_n692), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n580), .A2(new_n754), .A3(new_n678), .A4(new_n757), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT48), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n678), .A2(new_n757), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n660), .A2(new_n784), .A3(new_n383), .A4(new_n579), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n600), .A2(new_n608), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n578), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n692), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n708), .C1(new_n688), .C2(new_n690), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n580), .A3(new_n754), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n704), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n467), .A3(new_n647), .A4(new_n678), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT50), .Z(new_n794));
  NOR2_X1   g608(.A1(new_n600), .A2(new_n608), .ZN(new_n795));
  INV_X1    g609(.A(new_n703), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n785), .A2(new_n795), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n675), .A2(new_n676), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n774), .B1(new_n464), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n757), .A3(new_n791), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT51), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n783), .B(new_n792), .C1(new_n798), .C2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n321), .A2(new_n704), .A3(new_n632), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n679), .A2(new_n682), .A3(new_n805), .A4(new_n697), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n686), .B1(new_n790), .B2(new_n696), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT111), .A3(new_n679), .A4(new_n682), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n511), .A2(new_n620), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n627), .A2(new_n292), .A3(new_n596), .A4(new_n294), .ZN(new_n814));
  INV_X1    g628(.A(new_n632), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n597), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n626), .A2(new_n596), .A3(new_n594), .A4(new_n812), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n633), .A2(new_n819), .A3(KEYINPUT112), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n292), .A2(new_n627), .A3(new_n596), .A4(new_n294), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n383), .A2(new_n609), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n731), .A2(new_n590), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n818), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n618), .A2(new_n577), .A3(new_n640), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n758), .A2(new_n631), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n321), .A2(new_n826), .A3(new_n636), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n691), .A2(new_n648), .A3(new_n695), .A4(new_n732), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n744), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n811), .A2(new_n739), .A3(new_n740), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n649), .A2(new_n613), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n714), .A2(new_n716), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n641), .A2(KEYINPUT113), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n641), .A2(KEYINPUT113), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n631), .A2(new_n464), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n660), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n644), .B(new_n840), .C1(new_n667), .C2(new_n668), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n707), .A2(new_n711), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n832), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n644), .A2(new_n840), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n669), .A2(KEYINPUT52), .A3(new_n712), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n831), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n741), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n830), .A4(new_n811), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n832), .B1(new_n839), .B2(new_n660), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n669), .A2(new_n644), .A3(new_n712), .A4(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n843), .A2(new_n852), .A3(KEYINPUT114), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n843), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n847), .B(KEYINPUT54), .C1(new_n850), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT115), .B1(new_n824), .B2(new_n829), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT112), .B1(new_n633), .B2(new_n819), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n821), .A2(new_n822), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n591), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n744), .A2(new_n827), .A3(new_n828), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n820), .A4(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n383), .B(new_n718), .C1(new_n295), .C2(new_n320), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT103), .B1(new_n867), .B2(KEYINPUT42), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n735), .A2(new_n734), .A3(new_n719), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n868), .A2(new_n869), .B1(new_n780), .B2(new_n720), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(new_n806), .ZN(new_n871));
  INV_X1    g685(.A(new_n806), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n737), .A2(new_n872), .A3(KEYINPUT116), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n865), .B(new_n874), .C1(new_n853), .C2(new_n854), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n849), .B1(new_n831), .B2(new_n846), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n856), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n798), .A2(KEYINPUT117), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n794), .A2(new_n882), .A3(new_n797), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n883), .A3(new_n802), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n804), .B(new_n879), .C1(new_n880), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n692), .A2(new_n750), .A3(new_n464), .A4(new_n610), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n888), .A3(new_n647), .A4(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n885), .A2(new_n886), .B1(new_n660), .B2(new_n890), .ZN(G75));
  AOI21_X1  g705(.A(new_n302), .B1(new_n875), .B2(new_n876), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n498), .A2(new_n502), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n500), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n245), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(G51));
  AOI211_X1 g718(.A(new_n302), .B(new_n761), .C1(new_n875), .C2(new_n876), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n762), .B(KEYINPUT57), .Z(new_n906));
  AND3_X1   g720(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n671), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT119), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n875), .A2(new_n876), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n878), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n459), .B1(new_n915), .B2(new_n906), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n912), .B(new_n900), .C1(new_n916), .C2(new_n905), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  INV_X1    g733(.A(new_n541), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n900), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT120), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n899), .B1(new_n919), .B2(new_n920), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n925), .B(new_n926), .C1(new_n920), .C2(new_n919), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n879), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n606), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n606), .A2(new_n930), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n907), .B2(new_n908), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n933), .A2(new_n934), .A3(new_n900), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n900), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n879), .A2(new_n931), .B1(new_n604), .B2(new_n605), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT121), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n875), .B2(new_n876), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n899), .B1(new_n944), .B2(new_n629), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n365), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT122), .B1(new_n944), .B2(new_n629), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n582), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n245), .B1(new_n950), .B2(G224), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n811), .A2(new_n820), .A3(new_n861), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(new_n245), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n895), .B1(G898), .B2(new_n245), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n955), .B(new_n956), .Z(G69));
  NOR2_X1   g771(.A1(new_n269), .A2(new_n270), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n536), .B(KEYINPUT124), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n638), .B2(new_n245), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n767), .A2(new_n834), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n776), .B1(new_n780), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n669), .A2(new_n644), .A3(new_n712), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n770), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n848), .A2(new_n744), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n245), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n637), .A2(KEYINPUT125), .A3(new_n787), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n757), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT125), .B1(new_n637), .B2(new_n787), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n652), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n776), .B1(new_n731), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n965), .A2(new_n662), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n770), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n961), .B1(new_n980), .B2(new_n245), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n439), .B2(new_n638), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n961), .B2(KEYINPUT127), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n971), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n971), .B2(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n970), .B2(new_n953), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n990), .A2(new_n250), .A3(new_n311), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n954), .B2(new_n980), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n250), .A3(new_n311), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(new_n312), .B2(new_n655), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n847), .B(new_n994), .C1(new_n850), .C2(new_n855), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n900), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n991), .A2(new_n996), .ZN(G57));
endmodule


