//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(G57gat), .B(G85gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g014(.A(G120gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G113gat), .ZN(new_n217));
  INV_X1    g016(.A(G113gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G120gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n226), .A2(new_n228), .B1(KEYINPUT2), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT75), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n233), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n230), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  INV_X1    g044(.A(new_n229), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n236), .A2(KEYINPUT76), .A3(new_n229), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n224), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n227), .A2(G141gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n225), .A2(G148gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n242), .B1(new_n241), .B2(new_n233), .ZN(new_n256));
  AND4_X1   g055(.A1(new_n242), .A2(new_n232), .A3(new_n233), .A4(new_n236), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n215), .A2(new_n223), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n249), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT5), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n251), .B2(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT79), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n238), .A2(new_n243), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT76), .B1(new_n236), .B2(new_n229), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n270), .A2(new_n255), .B1(new_n272), .B2(new_n248), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT4), .B1(new_n273), .B2(new_n259), .ZN(new_n274));
  AND4_X1   g073(.A1(KEYINPUT4), .A2(new_n258), .A3(new_n249), .A4(new_n259), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n274), .A2(new_n275), .A3(new_n263), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT3), .B1(new_n244), .B2(new_n250), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n244), .C2(new_n250), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n249), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n224), .A4(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n266), .A2(new_n269), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n276), .A2(new_n268), .A3(new_n283), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT6), .B(new_n208), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n276), .A2(new_n268), .A3(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n207), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n289), .B2(new_n284), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n283), .A2(new_n291), .A3(new_n262), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n265), .B1(new_n264), .B2(KEYINPUT5), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n267), .A2(KEYINPUT79), .A3(new_n268), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n207), .B1(new_n295), .B2(new_n288), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n286), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(KEYINPUT22), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G211gat), .B(G218gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n316), .A2(KEYINPUT65), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT65), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n316), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n312), .B1(new_n324), .B2(new_n311), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT66), .B(KEYINPUT26), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n330), .B(KEYINPUT67), .C1(new_n331), .C2(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(new_n306), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n332), .A2(new_n333), .A3(new_n315), .A4(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n315), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n329), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(new_n334), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n333), .B1(new_n348), .B2(new_n332), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n326), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n351), .B(KEYINPUT71), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n332), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n315), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n338), .A3(new_n344), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n362), .B2(new_n326), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n363), .A2(KEYINPUT72), .A3(new_n354), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n305), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  AOI21_X1  g167(.A(new_n352), .B1(new_n350), .B2(new_n355), .ZN(new_n369));
  INV_X1    g168(.A(new_n354), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n362), .B2(new_n326), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n369), .A2(new_n371), .A3(new_n305), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT72), .B1(new_n363), .B2(new_n354), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n357), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n353), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n379), .B2(new_n305), .ZN(new_n380));
  INV_X1    g179(.A(new_n368), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(new_n375), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n297), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n351), .B1(new_n362), .B2(new_n326), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n350), .A2(new_n355), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n370), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n387), .B2(KEYINPUT72), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n304), .B1(new_n388), .B2(new_n378), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT73), .B1(new_n389), .B2(new_n372), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n391), .A3(new_n373), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n368), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n203), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n208), .B1(new_n284), .B2(new_n285), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n295), .A2(new_n288), .A3(new_n207), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n287), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(new_n286), .B1(new_n380), .B2(new_n382), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT73), .B(new_n372), .C1(new_n379), .C2(new_n305), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n365), .B2(new_n373), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n381), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n401), .A3(KEYINPUT80), .A4(new_n376), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  INV_X1    g205(.A(G50gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n304), .B(new_n355), .C1(new_n244), .C2(new_n250), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(G228gat), .A3(G233gat), .A4(new_n277), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n282), .A2(new_n355), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n304), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n282), .A2(KEYINPUT84), .A3(new_n355), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n417), .B(KEYINPUT83), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n281), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n304), .B2(new_n355), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n421), .A2(new_n273), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n304), .B1(new_n282), .B2(new_n355), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n419), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(G22gat), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n414), .A2(new_n415), .ZN(new_n427));
  INV_X1    g226(.A(new_n411), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G22gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n421), .A2(new_n273), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n418), .B1(new_n431), .B2(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n409), .B1(new_n434), .B2(KEYINPUT82), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436));
  AOI211_X1 g235(.A(new_n436), .B(new_n408), .C1(new_n426), .C2(new_n433), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n405), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n350), .A2(new_n224), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n362), .A2(new_n259), .A3(new_n326), .ZN(new_n440));
  INV_X1    g239(.A(G227gat), .ZN(new_n441));
  INV_X1    g240(.A(G233gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT34), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(KEYINPUT34), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n439), .B2(new_n440), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(KEYINPUT33), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(new_n456), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT69), .B(new_n449), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  INV_X1    g260(.A(new_n448), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT69), .A3(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n447), .B2(new_n448), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n457), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n416), .A2(new_n425), .A3(G22gat), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT82), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n408), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n434), .A2(KEYINPUT82), .A3(new_n409), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n404), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n438), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT35), .B1(new_n403), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n376), .A2(new_n383), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT85), .B1(new_n393), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n374), .A2(new_n375), .B1(new_n380), .B2(new_n382), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n401), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n397), .A2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n395), .A2(new_n396), .A3(new_n485), .A4(new_n287), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n286), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n475), .A2(new_n476), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n403), .C2(new_n474), .ZN(new_n491));
  AND4_X1   g290(.A1(new_n279), .A2(new_n280), .A3(new_n224), .A4(new_n282), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n274), .A2(new_n275), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n263), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT39), .C1(new_n263), .C2(new_n261), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n263), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n207), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT86), .B1(new_n497), .B2(new_n207), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT40), .B(new_n495), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n395), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n498), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT40), .B1(new_n504), .B2(new_n495), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n401), .A2(new_n479), .A3(new_n480), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n479), .B1(new_n401), .B2(new_n480), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n438), .A2(new_n473), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n368), .B1(new_n380), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n379), .A2(new_n304), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n369), .A2(new_n371), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n516), .B2(new_n305), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n374), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n487), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n512), .B1(new_n390), .B2(new_n392), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n514), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n511), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n482), .A2(new_n527), .A3(new_n506), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n467), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n460), .A2(new_n466), .A3(KEYINPUT70), .A4(KEYINPUT36), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n403), .B2(new_n511), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n490), .A2(new_n491), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n234), .ZN(new_n538));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n543), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n543), .B(new_n542), .C1(new_n546), .C2(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n554), .A2(G127gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(KEYINPUT94), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT16), .ZN(new_n558));
  AOI21_X1  g357(.A(G1gat), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  INV_X1    g360(.A(G8gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT95), .B(G8gat), .Z(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(KEYINPUT21), .B2(new_n551), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n554), .A2(G127gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n555), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n555), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n541), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n569), .A3(new_n540), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT15), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n576), .B2(new_n577), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT93), .B(G43gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n407), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n407), .A2(G43gat), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT15), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G29gat), .A2(G36gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR3_X1    g387(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n581), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n580), .A3(new_n591), .A4(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G99gat), .ZN(new_n602));
  INV_X1    g401(.A(G106gat), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT8), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n601), .B(new_n604), .C1(G85gat), .C2(G92gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT7), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR4_X1   g407(.A1(new_n608), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n610), .A2(KEYINPUT99), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(KEYINPUT99), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n612), .ZN(new_n618));
  INV_X1    g417(.A(new_n595), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n622), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n616), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n616), .B(new_n627), .C1(new_n621), .C2(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n629), .B1(KEYINPUT101), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n632), .B(KEYINPUT101), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n551), .A2(new_n613), .A3(new_n614), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(new_n644), .C1(new_n618), .C2(new_n551), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n551), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n644), .B1(new_n618), .B2(new_n551), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n640), .B1(new_n650), .B2(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n652), .B(new_n639), .C1(new_n647), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n575), .A2(new_n634), .A3(new_n636), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n565), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n597), .ZN(new_n657));
  NAND2_X1  g456(.A1(G229gat), .A2(G233gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n565), .A2(new_n619), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT18), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n565), .B(new_n619), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n658), .B(KEYINPUT13), .Z(new_n663));
  AOI22_X1  g462(.A1(new_n660), .A2(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n657), .A2(new_n659), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(KEYINPUT18), .A3(new_n658), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G113gat), .B(G141gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G197gat), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT11), .B(G169gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT12), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n660), .A2(new_n661), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(KEYINPUT96), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n667), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n655), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n202), .B1(new_n536), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n475), .A2(new_n476), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n483), .A2(new_n489), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n491), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n529), .A2(new_n535), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n297), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT104), .B(G1gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1324gat));
  INV_X1    g492(.A(new_n482), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n562), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n694), .B(new_n697), .C1(new_n682), .C2(new_n688), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT103), .B1(new_n687), .B2(new_n680), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n202), .B(new_n681), .C1(new_n685), .C2(new_n686), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n482), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n698), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n482), .B(new_n696), .C1(new_n699), .C2(new_n700), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n702), .B(new_n709), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1325gat));
  INV_X1    g510(.A(new_n689), .ZN(new_n712));
  INV_X1    g511(.A(new_n467), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n712), .A2(G15gat), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n534), .ZN(new_n715));
  OAI21_X1  g514(.A(G15gat), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n689), .A2(new_n511), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n634), .A2(new_n636), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n536), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n654), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n679), .A2(new_n575), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(G29gat), .A3(new_n297), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n687), .A2(new_n723), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n727), .B(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n297), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n728), .A2(G36gat), .A3(new_n694), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n738), .B2(new_n694), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(new_n582), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n728), .B2(new_n713), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n534), .A2(new_n582), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n738), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n750), .B(new_n746), .C1(new_n738), .C2(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1330gat));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n735), .A3(new_n511), .A4(new_n737), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT112), .B1(new_n725), .B2(new_n727), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n725), .A2(KEYINPUT112), .A3(new_n727), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n407), .A3(new_n511), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1331gat));
  NAND4_X1  g559(.A1(new_n679), .A2(new_n724), .A3(new_n575), .A4(new_n726), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n536), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n690), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n762), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n694), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n766), .B2(new_n715), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n762), .B2(new_n467), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n536), .A2(KEYINPUT114), .A3(new_n713), .A4(new_n761), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n772), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n773), .B1(new_n772), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1334gat));
  AND2_X1   g580(.A1(new_n438), .A2(new_n473), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(G78gat), .Z(G1335gat));
  INV_X1    g583(.A(new_n575), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n679), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT115), .Z(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n654), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n736), .A2(new_n690), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n733), .B2(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(new_n787), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n726), .A2(new_n599), .A3(new_n690), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n789), .A2(new_n599), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  NAND4_X1  g595(.A1(new_n732), .A2(new_n735), .A3(new_n482), .A4(new_n788), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n694), .A2(G92gat), .A3(new_n654), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n798), .B(new_n799), .C1(new_n794), .C2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n791), .A2(new_n793), .A3(new_n803), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(new_n800), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n798), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n802), .B1(new_n807), .B2(new_n799), .ZN(G1337gat));
  NAND4_X1  g607(.A1(new_n732), .A2(new_n735), .A3(new_n534), .A4(new_n788), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G99gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n726), .A2(new_n602), .A3(new_n467), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT117), .Z(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n794), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT118), .ZN(G1338gat));
  NAND4_X1  g613(.A1(new_n732), .A2(new_n735), .A3(new_n511), .A4(new_n788), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n782), .A2(G106gat), .A3(new_n654), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n816), .B(new_n817), .C1(new_n794), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n818), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n816), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(new_n817), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n655), .A2(new_n678), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n665), .A2(new_n658), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n662), .A2(new_n663), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n671), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n664), .A2(new_n666), .A3(new_n673), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n726), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n639), .B1(new_n647), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n647), .A2(new_n831), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n645), .A2(new_n642), .A3(new_n646), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n650), .A2(new_n639), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT55), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n724), .B(new_n830), .C1(new_n679), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n829), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n575), .B1(new_n842), .B2(new_n723), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n824), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n844), .A2(new_n297), .A3(new_n482), .A4(new_n511), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n467), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n218), .A3(new_n679), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n844), .A2(new_n297), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n483), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n678), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n851), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n850), .B2(new_n726), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n713), .A2(new_n216), .A3(new_n654), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n845), .B2(new_n854), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n846), .B2(new_n785), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n211), .A3(new_n575), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT119), .Z(G1342gat));
  NAND3_X1  g658(.A1(new_n850), .A2(new_n209), .A3(new_n723), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n846), .B2(new_n724), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n534), .A2(new_n782), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n694), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(G141gat), .A3(new_n679), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n534), .A2(new_n482), .A3(new_n297), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n723), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n785), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n827), .A2(new_n828), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n634), .B(new_n636), .C1(new_n872), .C2(new_n654), .ZN(new_n873));
  INV_X1    g672(.A(new_n840), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n678), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n871), .A2(new_n875), .B1(new_n655), .B2(new_n678), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n511), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n844), .A2(new_n878), .A3(new_n782), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n869), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n679), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n868), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(KEYINPUT120), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(new_n869), .C1(new_n877), .C2(new_n879), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n678), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT121), .B1(new_n887), .B2(G141gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n867), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n890), .B2(new_n882), .ZN(G1344gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  INV_X1    g691(.A(new_n866), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n892), .B(G148gat), .C1(new_n893), .C2(new_n726), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n878), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n877), .A2(new_n879), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(KEYINPUT122), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n726), .A3(new_n869), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n227), .B1(new_n899), .B2(KEYINPUT59), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n884), .A2(new_n886), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n892), .A3(new_n726), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  AOI21_X1  g702(.A(G155gat), .B1(new_n893), .B2(new_n575), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n575), .A2(G155gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT123), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n901), .B2(new_n906), .ZN(G1346gat));
  AOI21_X1  g706(.A(G162gat), .B1(new_n893), .B2(new_n723), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n724), .A2(new_n235), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n901), .B2(new_n909), .ZN(G1347gat));
  NOR4_X1   g709(.A1(new_n844), .A2(new_n690), .A3(new_n694), .A4(new_n474), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n678), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n726), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g714(.A(G183gat), .B1(new_n911), .B2(new_n575), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n575), .ZN(new_n918));
  OAI221_X1 g717(.A(new_n917), .B1(KEYINPUT124), .B2(KEYINPUT60), .C1(new_n339), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1350gat));
  NAND2_X1  g720(.A1(new_n911), .A2(new_n723), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G190gat), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n925), .ZN(new_n926));
  OAI221_X1 g725(.A(new_n926), .B1(KEYINPUT61), .B2(new_n925), .C1(G190gat), .C2(new_n922), .ZN(G1351gat));
  NAND4_X1  g726(.A1(new_n876), .A2(new_n297), .A3(new_n482), .A4(new_n865), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n678), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n694), .A2(new_n534), .A3(new_n690), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n898), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n678), .A2(G197gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n726), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G204gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n928), .A2(G204gat), .A3(new_n654), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n930), .A2(new_n299), .A3(new_n575), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n898), .A2(new_n575), .A3(new_n932), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n930), .B2(new_n723), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n723), .A2(G218gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n933), .B2(new_n948), .ZN(G1355gat));
endmodule


