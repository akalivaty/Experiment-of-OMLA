//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G29gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT15), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(KEYINPUT15), .B2(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(G1gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT16), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(G1gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n212), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n215), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n221), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n213), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n227), .B2(new_n213), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n222), .A2(KEYINPUT90), .A3(new_n211), .A4(new_n212), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n228), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n225), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n224), .A2(KEYINPUT18), .A3(new_n225), .A4(new_n228), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G169gat), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT12), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n237), .A3(new_n238), .A4(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G155gat), .ZN(new_n251));
  INV_X1    g050(.A(G162gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G141gat), .B(G148gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(KEYINPUT2), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G148gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(G141gat), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT76), .B(G148gat), .Z(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(G141gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n253), .B1(new_n262), .B2(new_n254), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  INV_X1    g067(.A(G113gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G120gat), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n274), .A2(KEYINPUT66), .A3(G127gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n272), .B2(KEYINPUT66), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n268), .B1(new_n266), .B2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g076(.A(G120gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G113gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n270), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n266), .A2(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n268), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n288), .B2(new_n276), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n265), .B(new_n273), .C1(new_n284), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT4), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n285), .A3(new_n276), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n273), .A4(new_n265), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(KEYINPUT77), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n290), .A2(new_n298), .A3(KEYINPUT4), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n264), .B(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n273), .B1(new_n284), .B2(new_n289), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n297), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n264), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n290), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n309), .B2(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n303), .A2(new_n304), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n307), .A2(new_n300), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n290), .B2(KEYINPUT4), .ZN(new_n315));
  INV_X1    g114(.A(new_n296), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n290), .A2(new_n314), .A3(KEYINPUT4), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n312), .B(new_n313), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT0), .ZN(new_n322));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n319), .A3(new_n324), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G169gat), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n332), .A2(KEYINPUT26), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT27), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT65), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n346));
  AOI21_X1  g145(.A(G190gat), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n344), .A2(new_n349), .A3(G190gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n339), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n355), .B2(new_n333), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  OR3_X1    g162(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n358), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n336), .B1(new_n332), .B2(new_n354), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT25), .A4(new_n353), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g174(.A1(G211gat), .A2(G218gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(KEYINPUT72), .B2(KEYINPUT22), .ZN(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n376), .A4(new_n378), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n373), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT75), .B1(new_n370), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT75), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n394), .B(new_n373), .C1(new_n351), .C2(new_n369), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n374), .B(new_n391), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n370), .A2(new_n392), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n351), .B2(new_n369), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n399), .B2(new_n391), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n374), .B(new_n400), .C1(new_n393), .C2(new_n395), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n396), .B2(new_n401), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n419), .C1(new_n420), .C2(new_n409), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n396), .A2(new_n401), .A3(new_n405), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n320), .A2(KEYINPUT6), .A3(new_n325), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n329), .A2(new_n418), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n422), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n417), .B2(KEYINPUT86), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT87), .A3(new_n329), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n402), .A2(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n412), .B1(new_n411), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n309), .B2(new_n301), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n308), .A2(KEYINPUT83), .A3(new_n290), .A4(new_n300), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT39), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n301), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT84), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n444), .A3(new_n301), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n324), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n324), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT84), .B(new_n442), .C1(new_n447), .C2(new_n440), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n422), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n446), .A2(new_n448), .A3(new_n326), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G228gat), .ZN(new_n454));
  INV_X1    g253(.A(G233gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n384), .B2(new_n387), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n380), .A2(new_n386), .A3(new_n382), .A4(new_n383), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT3), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n265), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n384), .A2(new_n385), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n386), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n302), .B(new_n257), .C1(new_n261), .C2(new_n263), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n463), .A2(new_n388), .B1(new_n371), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n457), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n371), .A3(new_n388), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n265), .B1(new_n467), .B2(new_n302), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n371), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n389), .B2(new_n390), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n456), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G22gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G50gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G22gat), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n466), .B(new_n478), .C1(new_n468), .C2(new_n471), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n468), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n384), .A2(new_n387), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n371), .A3(new_n459), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n302), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n264), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n456), .B1(new_n486), .B2(new_n470), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n481), .B(G22gat), .C1(new_n482), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n479), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n472), .B2(G22gat), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT81), .B(new_n476), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n302), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n264), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n465), .A2(new_n457), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n470), .B1(new_n265), .B2(new_n460), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n494), .A2(new_n495), .B1(new_n496), .B2(new_n457), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT80), .B1(new_n497), .B2(new_n478), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n488), .A3(new_n479), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT81), .B1(new_n499), .B2(new_n476), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n480), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n453), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n434), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n476), .B1(new_n489), .B2(new_n490), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n491), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n508), .B2(new_n480), .ZN(new_n509));
  INV_X1    g308(.A(new_n480), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT82), .B(new_n510), .C1(new_n507), .C2(new_n491), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n452), .B1(new_n329), .B2(new_n424), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n351), .A2(new_n369), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n304), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n370), .A2(new_n294), .A3(new_n273), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT33), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n521), .B2(KEYINPUT32), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT34), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n521), .B(KEYINPUT32), .C1(new_n522), .C2(new_n529), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n531), .B2(new_n537), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT71), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n516), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT36), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n503), .A2(new_n515), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(KEYINPUT88), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n538), .B2(new_n540), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n514), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n501), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n513), .A2(new_n501), .A3(new_n543), .A4(new_n541), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n250), .B1(new_n547), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(G57gat), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT9), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n561), .B2(G57gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT92), .B1(new_n563), .B2(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n561), .A3(G57gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n563), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n566), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT93), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT95), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n584), .A2(new_n586), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n560), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  INV_X1    g390(.A(new_n560), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n587), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n222), .B1(new_n582), .B2(new_n581), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n590), .A2(new_n593), .A3(new_n600), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT8), .ZN(new_n609));
  OAI22_X1  g408(.A1(new_n606), .A2(new_n609), .B1(G85gat), .B2(G92gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  OR2_X1    g410(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n612));
  AND3_X1   g411(.A1(KEYINPUT96), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT97), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n611), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(KEYINPUT96), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n608), .B(new_n610), .C1(new_n615), .C2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n608), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(new_n610), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n215), .B(new_n223), .C1(new_n622), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n622), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n628), .A2(new_n213), .B1(KEYINPUT41), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n605), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n630), .A3(new_n605), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(new_n631), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n602), .A2(new_n603), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n625), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n608), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n570), .A2(new_n580), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n624), .A2(new_n623), .A3(new_n625), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n581), .B1(new_n626), .B2(new_n622), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n649), .A2(new_n650), .A3(new_n654), .A4(new_n651), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n644), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n649), .A2(new_n650), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n643), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G120gat), .B(G148gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n658), .A2(new_n660), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n559), .A2(new_n641), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n329), .A2(new_n424), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n217), .ZN(G1324gat));
  INV_X1    g473(.A(new_n671), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n452), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n677), .A2(KEYINPUT101), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n226), .B1(new_n675), .B2(new_n452), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n677), .B1(new_n683), .B2(new_n678), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n679), .B1(new_n682), .B2(new_n684), .ZN(G1325gat));
  NOR3_X1   g484(.A1(new_n544), .A2(KEYINPUT102), .A3(new_n545), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n540), .A2(new_n539), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n548), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n540), .A2(new_n539), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT36), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n545), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n671), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n549), .A2(new_n552), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(G15gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n671), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n510), .B1(new_n507), .B2(new_n491), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n504), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n671), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n547), .A2(new_n558), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n640), .A2(new_n637), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n602), .A2(new_n603), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n710), .A3(new_n669), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n249), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n672), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n203), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n554), .A2(new_n501), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n434), .A2(new_n502), .B1(new_n512), .B2(new_n514), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n694), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(new_n709), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n709), .A2(new_n717), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n710), .B1(new_n707), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n250), .A2(new_n669), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n714), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G29gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n727), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n451), .A2(G36gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT103), .B1(new_n712), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n559), .A2(new_n733), .A3(new_n711), .A4(new_n729), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n731), .A2(KEYINPUT105), .A3(new_n732), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n452), .A3(new_n725), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G36gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n731), .A2(new_n734), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT104), .B1(new_n742), .B2(KEYINPUT46), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n739), .B(new_n741), .C1(new_n743), .C2(new_n744), .ZN(G1329gat));
  OAI21_X1  g544(.A(KEYINPUT102), .B1(new_n544), .B2(new_n545), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n691), .A2(new_n687), .A3(new_n692), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n721), .A2(new_n723), .A3(new_n748), .A4(new_n725), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G43gat), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n712), .A2(G43gat), .A3(new_n697), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1330gat));
  NAND4_X1  g553(.A1(new_n721), .A2(new_n723), .A3(new_n512), .A4(new_n725), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n703), .A2(G50gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n712), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT48), .B1(new_n757), .B2(new_n760), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n721), .A2(new_n723), .A3(new_n701), .A4(new_n725), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(G50gat), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n762), .A2(KEYINPUT48), .B1(new_n763), .B2(new_n765), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n670), .A2(new_n249), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n641), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT107), .Z(new_n769));
  OAI21_X1  g568(.A(KEYINPUT108), .B1(new_n720), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n503), .A2(new_n515), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n558), .B1(new_n771), .B2(new_n748), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n773));
  INV_X1    g572(.A(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n672), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n563), .ZN(G1332gat));
  XNOR2_X1  g577(.A(new_n451), .B(KEYINPUT109), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n770), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n561), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n783), .A2(new_n786), .A3(new_n561), .A4(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1333gat));
  OAI21_X1  g589(.A(new_n567), .B1(new_n776), .B2(new_n697), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n770), .A2(new_n775), .A3(G71gat), .A4(new_n748), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g593(.A1(new_n776), .A2(new_n703), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n568), .ZN(G1335gat));
  NAND2_X1  g595(.A1(new_n724), .A2(new_n767), .ZN(new_n797));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797), .B2(new_n672), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n249), .B(new_n710), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n772), .A2(new_n708), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n803), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n772), .A2(new_n708), .A3(new_n805), .A4(new_n801), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n672), .A2(G85gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n669), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n798), .A2(new_n809), .ZN(G1336gat));
  INV_X1    g609(.A(G92gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n779), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n721), .A2(new_n723), .A3(new_n767), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(KEYINPUT114), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n724), .A2(new_n815), .A3(new_n767), .A4(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n779), .A2(G92gat), .A3(new_n670), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n807), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n721), .A2(new_n723), .A3(new_n452), .A4(new_n767), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G92gat), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n818), .B(KEYINPUT113), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n806), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(G1337gat));
  OAI21_X1  g626(.A(G99gat), .B1(new_n797), .B2(new_n694), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n697), .A2(G99gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n669), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1338gat));
  NOR3_X1   g630(.A1(new_n501), .A2(G106gat), .A3(new_n670), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT115), .Z(new_n833));
  NAND2_X1  g632(.A1(new_n807), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n721), .A2(new_n723), .A3(new_n701), .A4(new_n767), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(G106gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n721), .A2(new_n723), .A3(new_n512), .A4(new_n767), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G106gat), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n804), .A2(KEYINPUT116), .A3(new_n806), .A4(new_n833), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n836), .B2(new_n843), .ZN(G1339gat));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n643), .A3(new_n655), .A4(new_n656), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n666), .B1(new_n658), .B2(KEYINPUT54), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n655), .A2(new_n656), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n643), .B1(new_n851), .B2(new_n846), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n665), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n850), .A2(new_n249), .A3(new_n856), .A4(new_n668), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n235), .A2(new_n236), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n225), .B1(new_n224), .B2(new_n228), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n244), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n248), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n708), .B1(new_n669), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n850), .A2(new_n668), .A3(new_n856), .A4(new_n861), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n708), .ZN(new_n865));
  INV_X1    g664(.A(new_n710), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n641), .A2(new_n250), .A3(new_n670), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n703), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT117), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n812), .A2(new_n672), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n696), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n269), .A3(new_n250), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n710), .B1(new_n864), .B2(new_n708), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n868), .B1(new_n876), .B2(new_n863), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n672), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n701), .A2(new_n689), .A3(new_n690), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n812), .ZN(new_n881));
  AOI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n249), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n875), .A2(new_n882), .ZN(G1340gat));
  OAI21_X1  g682(.A(G120gat), .B1(new_n874), .B2(new_n670), .ZN(new_n884));
  INV_X1    g683(.A(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n669), .A2(new_n278), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT118), .Z(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n874), .B2(new_n866), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n885), .A2(G127gat), .A3(new_n866), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1342gat));
  OAI21_X1  g690(.A(G134gat), .B1(new_n874), .B2(new_n709), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n452), .A2(new_n709), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n274), .A3(new_n879), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT56), .Z(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1343gat));
  NAND3_X1  g695(.A1(new_n746), .A2(new_n873), .A3(new_n747), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n877), .A2(new_n703), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n870), .A2(KEYINPUT57), .A3(new_n512), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n877), .B2(new_n501), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT119), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n249), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G141gat), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n748), .A2(new_n501), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(new_n878), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n779), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n250), .A2(G141gat), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n906), .B(new_n907), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n909), .A2(new_n779), .A3(new_n911), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n902), .A2(KEYINPUT119), .A3(new_n903), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n870), .A2(new_n900), .A3(new_n512), .A4(KEYINPUT57), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n694), .A3(new_n873), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT120), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n919), .A3(new_n904), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n249), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n914), .B1(new_n921), .B2(G141gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n913), .B1(new_n922), .B2(new_n907), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT121), .B(new_n913), .C1(new_n922), .C2(new_n907), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1344gat));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n918), .A2(new_n920), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n670), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n930), .B2(new_n260), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n669), .A2(new_n260), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n877), .A2(new_n703), .A3(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n898), .B1(new_n870), .B2(new_n701), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(new_n670), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n897), .A2(KEYINPUT122), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n897), .A2(KEYINPUT122), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n939));
  OAI221_X1 g738(.A(new_n931), .B1(new_n910), .B2(new_n932), .C1(new_n938), .C2(new_n939), .ZN(G1345gat));
  INV_X1    g739(.A(new_n929), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n710), .A2(G155gat), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT123), .Z(new_n943));
  NAND3_X1  g742(.A1(new_n909), .A2(new_n710), .A3(new_n779), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n941), .A2(new_n943), .B1(new_n251), .B2(new_n944), .ZN(G1346gat));
  NAND3_X1  g744(.A1(new_n909), .A2(new_n252), .A3(new_n893), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  OAI21_X1  g746(.A(G162gat), .B1(new_n929), .B2(new_n709), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n672), .A2(new_n452), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n697), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n872), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n330), .A3(new_n250), .ZN(new_n953));
  AND4_X1   g752(.A1(new_n672), .A2(new_n870), .A3(new_n879), .A4(new_n812), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n249), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n955), .ZN(G1348gat));
  OAI21_X1  g755(.A(G176gat), .B1(new_n952), .B2(new_n670), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n331), .A3(new_n669), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n952), .B2(new_n866), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT60), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n954), .A2(new_n341), .A3(new_n343), .A4(new_n710), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n960), .B(new_n962), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n961), .A2(KEYINPUT60), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n359), .A3(new_n708), .ZN(new_n970));
  OAI21_X1  g769(.A(G190gat), .B1(new_n952), .B2(new_n709), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n877), .A2(new_n714), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n908), .A2(new_n812), .A3(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n249), .ZN(new_n978));
  NOR4_X1   g777(.A1(new_n933), .A2(new_n934), .A3(new_n748), .A4(new_n950), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n249), .A2(G197gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NAND4_X1  g780(.A1(new_n935), .A2(new_n672), .A3(new_n452), .A4(new_n694), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  OR3_X1    g782(.A1(new_n976), .A2(G204gat), .A3(new_n670), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n983), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(G1353gat));
  OR3_X1    g788(.A1(new_n976), .A2(G211gat), .A3(new_n866), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n979), .A2(new_n710), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  INV_X1    g793(.A(G218gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n977), .A2(new_n995), .A3(new_n708), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n979), .A2(new_n708), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n997), .B2(new_n995), .ZN(G1355gat));
endmodule


