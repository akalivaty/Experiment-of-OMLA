//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT64), .B1(new_n187), .B2(G134), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(G134), .B2(new_n187), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n190), .A2(KEYINPUT11), .A3(G137), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n195), .B(new_n196), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n204), .A2(KEYINPUT1), .A3(G146), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT65), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n202), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n201), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n204), .A2(G146), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n209), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT0), .A4(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n226), .B2(new_n200), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT30), .B1(new_n218), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n224), .ZN(new_n229));
  INV_X1    g043(.A(new_n200), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n192), .A2(KEYINPUT11), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n197), .A2(new_n187), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n195), .B1(new_n233), .B2(new_n196), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n229), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  INV_X1    g050(.A(new_n217), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n208), .B2(new_n213), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n235), .B(new_n236), .C1(new_n238), .C2(new_n201), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G113), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G116), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n242), .B(new_n244), .C1(new_n246), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n244), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n240), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n215), .B1(new_n221), .B2(new_n209), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n211), .B1(new_n255), .B2(new_n210), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n217), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n201), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n265), .A3(new_n235), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n254), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n218), .A2(new_n264), .A3(new_n227), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n240), .B2(new_n253), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT31), .A3(new_n272), .ZN(new_n278));
  INV_X1    g092(.A(new_n253), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n260), .B2(new_n235), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n280), .B2(new_n276), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n266), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT67), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n272), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n275), .A2(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT32), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n287), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT31), .B1(new_n277), .B2(new_n272), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n279), .B1(new_n228), .B2(new_n239), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n294), .A2(new_n274), .A3(new_n276), .A4(new_n287), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n289), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n281), .A2(new_n285), .A3(new_n284), .A4(new_n272), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n287), .B1(new_n294), .B2(new_n276), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n304), .A3(new_n300), .A4(new_n301), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n265), .B1(new_n260), .B2(new_n235), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT28), .B1(new_n306), .B2(new_n276), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n287), .A2(new_n300), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n284), .A3(new_n285), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n303), .A2(new_n305), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n291), .A2(new_n298), .B1(new_n313), .B2(G472), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G137), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(KEYINPUT69), .A3(G125), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n202), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI211_X1 g145(.A(KEYINPUT70), .B(new_n202), .C1(new_n326), .C2(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n247), .B2(G128), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(new_n335), .C1(G119), .C2(new_n215), .ZN(new_n336));
  XNOR2_X1  g150(.A(G119), .B(G128), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT24), .B(G110), .Z(new_n338));
  OAI22_X1  g152(.A1(new_n336), .A2(G110), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n320), .A2(new_n322), .A3(new_n202), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n331), .A2(new_n332), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(G110), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n326), .A2(new_n328), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n326), .A2(new_n202), .A3(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n318), .B1(new_n342), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n329), .A2(new_n330), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(new_n340), .A3(new_n352), .A4(new_n339), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n317), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n355), .A3(new_n310), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n350), .A2(new_n355), .A3(KEYINPUT25), .A4(new_n310), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G217), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G234), .B2(new_n310), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n362), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n350), .A2(new_n355), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n362), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT72), .B1(new_n314), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n303), .A2(new_n305), .A3(new_n312), .ZN(new_n372));
  INV_X1    g186(.A(G472), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n296), .A2(new_n297), .A3(new_n289), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n297), .B1(new_n296), .B2(new_n289), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n245), .A2(G122), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT86), .A2(G122), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT86), .A2(G122), .ZN(new_n388));
  OAI21_X1  g202(.A(G116), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n382), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n215), .A2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n204), .A2(G128), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n204), .A2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n215), .A2(G143), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n190), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n382), .A3(new_n383), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n381), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n383), .B(KEYINPUT14), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n245), .B1(new_n404), .B2(new_n386), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(KEYINPUT90), .A3(new_n398), .A4(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n383), .ZN(new_n409));
  OAI21_X1  g223(.A(G107), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n398), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT13), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n412), .B(new_n394), .C1(new_n392), .C2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n391), .B1(KEYINPUT13), .B2(new_n395), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT87), .B1(new_n394), .B2(new_n413), .ZN(new_n416));
  OAI211_X1 g230(.A(G134), .B(new_n414), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n396), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT88), .A4(new_n190), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n411), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n410), .A2(new_n398), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT89), .B1(new_n425), .B2(new_n417), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n408), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n428), .A2(new_n361), .A3(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n423), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(KEYINPUT89), .A3(new_n417), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n431), .A2(new_n432), .B1(new_n400), .B2(new_n407), .ZN(new_n433));
  INV_X1    g247(.A(new_n429), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n435), .A3(new_n310), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(G952), .A3(new_n268), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n436), .A2(new_n438), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n439), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT81), .B(G143), .ZN(new_n451));
  INV_X1    g265(.A(G214), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(G237), .A3(G953), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n267), .A2(new_n268), .A3(G214), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(KEYINPUT81), .B2(new_n204), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT17), .B(G131), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n347), .A2(new_n348), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n347), .A2(new_n460), .A3(new_n348), .A4(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(G131), .B1(new_n454), .B2(new_n456), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n453), .B1(new_n464), .B2(G143), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n195), .C1(new_n453), .C2(new_n451), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n459), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n324), .A2(new_n325), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G146), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n340), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT82), .A2(KEYINPUT18), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(G131), .B(new_n474), .C1(new_n454), .C2(new_n456), .ZN(new_n475));
  OAI221_X1 g289(.A(new_n465), .B1(new_n195), .B2(new_n473), .C1(new_n453), .C2(new_n451), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G113), .B(G122), .ZN(new_n478));
  INV_X1    g292(.A(G104), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT83), .Z(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n477), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n467), .B1(new_n458), .B2(KEYINPUT84), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n461), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT85), .A3(new_n481), .ZN(new_n488));
  INV_X1    g302(.A(new_n487), .ZN(new_n489));
  INV_X1    g303(.A(new_n480), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n484), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G475), .B1(new_n491), .B2(G902), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n320), .A2(new_n322), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n470), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n202), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n462), .A2(new_n466), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n351), .A2(new_n498), .A3(new_n499), .A4(new_n352), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n480), .B1(new_n500), .B2(new_n477), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n482), .A2(new_n483), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT85), .B1(new_n487), .B2(new_n481), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G475), .A2(G902), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n493), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n501), .B1(new_n484), .B2(new_n488), .ZN(new_n508));
  INV_X1    g322(.A(new_n506), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n508), .A2(KEYINPUT20), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n450), .B(new_n492), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n513));
  OAI21_X1  g327(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT3), .B1(new_n479), .B2(G107), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT3), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n382), .A3(G104), .ZN(new_n519));
  INV_X1    g333(.A(G101), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n479), .A2(G107), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n382), .A2(G104), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n521), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(G101), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT73), .B(new_n520), .C1(new_n524), .C2(new_n521), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n238), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G104), .B(G107), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT73), .B1(new_n530), .B2(new_n520), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n523), .A3(G101), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n217), .A2(new_n255), .A3(new_n210), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n522), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n226), .A2(new_n200), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT12), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n536), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n533), .A2(new_n545), .A3(new_n522), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n544), .A2(new_n258), .A3(KEYINPUT10), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT10), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(G101), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(G101), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n229), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n226), .A2(new_n557), .A3(new_n200), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(new_n549), .A3(new_n555), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G140), .ZN(new_n561));
  INV_X1    g375(.A(G227), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G953), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n561), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AND4_X1   g379(.A1(new_n541), .A2(new_n543), .A3(new_n560), .A4(new_n565), .ZN(new_n566));
  AND4_X1   g380(.A1(KEYINPUT10), .A2(new_n544), .A3(new_n258), .A4(new_n546), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n549), .A2(new_n555), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n537), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n569), .B2(new_n560), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n516), .B(new_n310), .C1(new_n566), .C2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n560), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n550), .B(new_n553), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(new_n229), .B1(new_n548), .B2(new_n535), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n538), .B1(new_n576), .B2(new_n547), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n564), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n541), .A2(new_n543), .A3(new_n560), .A4(new_n565), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT78), .A3(new_n516), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n560), .A2(new_n565), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n577), .B1(new_n583), .B2(KEYINPUT77), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n560), .A2(new_n585), .A3(new_n565), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n541), .A2(new_n543), .A3(new_n560), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n584), .A2(new_n586), .B1(new_n587), .B2(new_n564), .ZN(new_n588));
  OAI21_X1  g402(.A(G469), .B1(new_n588), .B2(G902), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n515), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G210), .B1(G237), .B2(G902), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT80), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n224), .A2(G125), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n258), .B2(G125), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(G224), .A3(new_n268), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n268), .A2(G224), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(new_n594), .C1(new_n258), .C2(G125), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n252), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n247), .A2(G116), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT5), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n241), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n544), .A2(new_n546), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n552), .A2(new_n554), .A3(new_n253), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n608), .ZN(new_n612));
  XNOR2_X1  g426(.A(G110), .B(G122), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT6), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n613), .B1(new_n609), .B2(new_n610), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT6), .A3(new_n612), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n600), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT7), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n597), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n599), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n595), .A2(new_n622), .A3(new_n597), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n606), .A2(new_n528), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n613), .B(KEYINPUT8), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n606), .A2(new_n528), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n616), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n593), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n620), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n619), .A2(new_n612), .B1(KEYINPUT6), .B2(new_n616), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n599), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n592), .A3(new_n631), .ZN(new_n637));
  OAI21_X1  g451(.A(G214), .B1(G237), .B2(G902), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n512), .A2(new_n513), .A3(new_n590), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n590), .A2(new_n639), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT92), .B1(new_n641), .B2(new_n511), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n380), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n505), .A2(new_n493), .A3(new_n506), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT20), .B1(new_n508), .B2(new_n509), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n489), .A2(new_n490), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n503), .B2(new_n504), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n310), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n646), .A2(new_n647), .B1(new_n650), .B2(G475), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n436), .A2(new_n437), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n429), .B1(new_n433), .B2(KEYINPUT94), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT94), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n427), .A2(new_n655), .A3(new_n434), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n656), .A3(KEYINPUT33), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT95), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n654), .A2(new_n656), .A3(new_n659), .A4(KEYINPUT33), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n430), .A2(new_n435), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n662));
  AOI22_X1  g476(.A1(new_n658), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n437), .A2(G902), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n653), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n645), .B1(new_n651), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n492), .B1(new_n507), .B2(new_n510), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n658), .A2(new_n660), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n661), .A2(new_n662), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n652), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n667), .A2(KEYINPUT96), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n296), .A2(new_n310), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G472), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n290), .B2(new_n288), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n447), .A3(new_n370), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n590), .A2(new_n639), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  NAND2_X1  g495(.A1(new_n439), .A2(new_n449), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n667), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n677), .A2(new_n678), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n353), .A2(new_n354), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n318), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n368), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n365), .A2(new_n366), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n642), .A2(new_n640), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  NAND3_X1  g510(.A1(new_n365), .A2(new_n366), .A3(new_n691), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n376), .A2(new_n590), .A3(new_n639), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n442), .B(KEYINPUT97), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(G900), .B2(new_n443), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT98), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n314), .A2(new_n692), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n704));
  INV_X1    g518(.A(new_n700), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n667), .A2(new_n683), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n678), .A2(new_n703), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  NOR2_X1   g523(.A1(new_n571), .A2(new_n572), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT78), .B1(new_n580), .B2(new_n516), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n589), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n514), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n700), .B(KEYINPUT39), .Z(new_n714));
  OR2_X1    g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n633), .A2(new_n637), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n374), .A2(new_n375), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n306), .A2(new_n276), .ZN(new_n722));
  AOI21_X1  g536(.A(G902), .B1(new_n722), .B2(new_n287), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n272), .B1(new_n294), .B2(new_n276), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n373), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n728));
  INV_X1    g542(.A(new_n638), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n651), .A2(new_n697), .A3(new_n683), .A4(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n716), .A2(new_n727), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  NOR3_X1   g546(.A1(new_n651), .A2(new_n665), .A3(new_n705), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n678), .A2(new_n703), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NOR2_X1   g549(.A1(new_n580), .A2(new_n516), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AND4_X1   g551(.A1(KEYINPUT100), .A2(new_n582), .A3(new_n514), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n573), .B2(new_n581), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT100), .B1(new_n739), .B2(new_n514), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n291), .A2(new_n298), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n313), .A2(G472), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n370), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n633), .A2(new_n637), .A3(new_n448), .A4(new_n638), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n673), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND2_X1  g563(.A1(new_n651), .A2(new_n682), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n745), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n514), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n739), .A2(KEYINPUT100), .A3(new_n514), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n744), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NOR3_X1   g571(.A1(new_n314), .A2(new_n511), .A3(new_n692), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n741), .A2(new_n758), .A3(new_n639), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND4_X1  g574(.A1(new_n633), .A2(new_n637), .A3(new_n682), .A4(new_n638), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n651), .A3(new_n447), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT102), .B(G472), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n674), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT101), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n307), .A2(new_n284), .A3(new_n285), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n275), .A2(new_n278), .B1(new_n287), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n767), .B2(new_n290), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n287), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n293), .B2(new_n295), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT101), .A3(new_n289), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n370), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n762), .A2(new_n773), .A3(new_n754), .A4(new_n755), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND3_X1  g589(.A1(new_n667), .A2(new_n671), .A3(new_n700), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n692), .A3(new_n772), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n639), .A3(new_n741), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  AOI21_X1  g593(.A(new_n311), .B1(new_n302), .B2(KEYINPUT68), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n373), .B1(new_n780), .B2(new_n305), .ZN(new_n781));
  OAI211_X1 g595(.A(KEYINPUT42), .B(new_n378), .C1(new_n721), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n776), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n729), .B1(new_n633), .B2(new_n637), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT103), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n515), .B1(new_n712), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n582), .A2(KEYINPUT103), .A3(new_n589), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n783), .A2(new_n784), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n717), .A2(new_n638), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n786), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n785), .A2(KEYINPUT104), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n789), .A3(new_n795), .A4(new_n790), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n744), .A2(new_n733), .A3(KEYINPUT42), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT105), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n787), .A3(new_n744), .A4(new_n733), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n792), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n195), .ZN(G33));
  NAND4_X1  g616(.A1(new_n791), .A2(new_n787), .A3(new_n744), .A4(new_n706), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G134), .ZN(G36));
  NAND2_X1  g618(.A1(new_n794), .A2(new_n795), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n667), .A2(new_n665), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT43), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n676), .A2(new_n697), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT44), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT107), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(G469), .B1(new_n588), .B2(KEYINPUT45), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT106), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n814), .A2(KEYINPUT106), .B1(KEYINPUT45), .B2(new_n588), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(G469), .A2(G902), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n582), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n514), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n714), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n813), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT107), .B1(new_n811), .B2(new_n812), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(new_n187), .ZN(G39));
  XOR2_X1   g643(.A(new_n824), .B(KEYINPUT47), .Z(new_n830));
  NOR3_X1   g644(.A1(new_n805), .A2(new_n376), .A3(new_n378), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n733), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G140), .ZN(G42));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  INV_X1    g648(.A(new_n699), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n807), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n370), .A3(new_n772), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n805), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n841));
  INV_X1    g655(.A(new_n739), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n514), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n830), .B2(KEYINPUT112), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n754), .A2(new_n755), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n719), .A3(new_n638), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n847), .A2(new_n837), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n837), .A2(new_n850), .B1(new_n847), .B2(new_n848), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(new_n847), .B2(new_n848), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n805), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n726), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n858), .A2(new_n442), .A3(new_n370), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(KEYINPUT117), .A3(new_n860), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n651), .A3(new_n665), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n772), .A2(new_n692), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  INV_X1    g681(.A(new_n836), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n857), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g683(.A(KEYINPUT116), .B(new_n836), .C1(new_n855), .C2(new_n856), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n853), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n834), .B1(new_n846), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n837), .A2(new_n639), .A3(new_n741), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(G952), .A3(new_n268), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n863), .A2(new_n864), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n673), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n744), .B1(new_n869), .B2(new_n870), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT48), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n839), .B1(new_n830), .B2(new_n843), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT51), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n873), .B(new_n882), .C1(new_n872), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n792), .A2(new_n798), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n799), .A2(new_n800), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n747), .A2(new_n759), .A3(new_n756), .A4(new_n774), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n791), .A2(new_n777), .A3(new_n787), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n667), .A2(new_n682), .A3(new_n705), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n787), .A2(new_n590), .A3(new_n703), .A4(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n803), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n677), .A2(new_n678), .A3(new_n667), .A4(new_n671), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n643), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n694), .A2(new_n685), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n694), .A2(new_n901), .A3(new_n685), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n708), .A2(new_n778), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT109), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT109), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n708), .A2(new_n907), .A3(new_n778), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n712), .A2(new_n788), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n365), .A2(new_n366), .A3(new_n691), .A4(new_n700), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n514), .A3(new_n790), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n789), .A2(KEYINPUT110), .A3(new_n790), .A4(new_n910), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n639), .A2(new_n667), .A3(new_n682), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n726), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n917), .A2(KEYINPUT52), .A3(new_n734), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n906), .A2(new_n908), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n708), .A2(new_n734), .A3(new_n778), .A4(new_n917), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT52), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n904), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n920), .B(KEYINPUT52), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n889), .B1(new_n886), .B2(new_n887), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n901), .B1(new_n694), .B2(new_n685), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n897), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(new_n929), .A3(new_n902), .A4(new_n894), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT53), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n931), .A3(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n894), .A2(KEYINPUT53), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n903), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT111), .B1(new_n801), .B2(new_n889), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT111), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n888), .A2(new_n936), .A3(new_n890), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n923), .A2(new_n934), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n924), .B1(new_n926), .B2(new_n930), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n885), .A2(new_n942), .B1(G952), .B2(G953), .ZN(new_n943));
  NOR4_X1   g757(.A1(new_n858), .A2(new_n515), .A3(new_n729), .A4(new_n370), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n719), .B1(KEYINPUT49), .B2(new_n842), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n842), .A2(KEYINPUT49), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n806), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(G75));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n950));
  INV_X1    g764(.A(new_n933), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n937), .A3(new_n951), .A4(new_n935), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n708), .A2(new_n907), .A3(new_n778), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n907), .B1(new_n708), .B2(new_n778), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g769(.A1(new_n955), .A2(new_n918), .B1(new_n921), .B2(new_n920), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n920), .B(new_n921), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n904), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(G902), .B(new_n592), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n634), .A2(new_n635), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n600), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n636), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT55), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n949), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  AOI211_X1 g782(.A(KEYINPUT118), .B(new_n968), .C1(new_n960), .C2(new_n961), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n310), .B1(new_n938), .B2(new_n939), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT119), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n592), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n961), .A3(new_n968), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n268), .A2(G952), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n970), .A2(new_n978), .ZN(G51));
  INV_X1    g793(.A(KEYINPUT120), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n310), .B(new_n817), .C1(new_n938), .C2(new_n939), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n818), .B(KEYINPUT57), .Z(new_n982));
  AND3_X1   g796(.A1(new_n938), .A2(new_n940), .A3(new_n939), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n578), .A2(new_n579), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n980), .B1(new_n987), .B2(new_n976), .ZN(new_n988));
  INV_X1    g802(.A(new_n986), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT54), .B1(new_n957), .B2(new_n959), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n941), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n991), .B2(new_n982), .ZN(new_n992));
  OAI211_X1 g806(.A(KEYINPUT120), .B(new_n977), .C1(new_n992), .C2(new_n981), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(new_n993), .ZN(G54));
  NAND3_X1  g808(.A1(new_n972), .A2(KEYINPUT58), .A3(G475), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n995), .A2(KEYINPUT121), .A3(new_n508), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n977), .B1(new_n995), .B2(new_n508), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT121), .B1(new_n995), .B2(new_n508), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(G60));
  NAND2_X1  g813(.A1(G478), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT59), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n663), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n990), .B2(new_n941), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT122), .B1(new_n1005), .B2(new_n977), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT122), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1004), .A2(new_n1007), .A3(new_n976), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n663), .B1(new_n942), .B2(new_n1002), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(G63));
  NAND2_X1  g824(.A1(G217), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT123), .Z(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT60), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n938), .B2(new_n939), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n690), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1015), .B(new_n977), .C1(new_n367), .C2(new_n1014), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G66));
  INV_X1    g832(.A(G224), .ZN(new_n1019));
  OAI21_X1  g833(.A(G953), .B1(new_n445), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n903), .A2(new_n889), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n963), .B1(G898), .B2(new_n268), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(G69));
  XOR2_X1   g838(.A(new_n497), .B(KEYINPUT124), .Z(new_n1025));
  XNOR2_X1  g839(.A(new_n240), .B(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  OAI211_X1 g841(.A(G900), .B(G953), .C1(new_n1027), .C2(G227), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(G227), .B2(new_n1027), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n888), .A2(new_n803), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n915), .A2(new_n314), .A3(new_n370), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n825), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n832), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n828), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n955), .A2(new_n734), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1033), .A2(KEYINPUT127), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1034), .A2(new_n832), .A3(new_n1035), .A4(new_n1032), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT127), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(G953), .B1(new_n1040), .B2(new_n1027), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1035), .A2(new_n731), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT62), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1035), .A2(KEYINPUT62), .A3(new_n731), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n684), .B1(new_n667), .B2(new_n671), .ZN(new_n1047));
  OR3_X1    g861(.A1(new_n1047), .A2(new_n715), .A3(new_n805), .ZN(new_n1048));
  INV_X1    g862(.A(new_n380), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(KEYINPUT125), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1051), .B1(new_n826), .B2(new_n827), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT126), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n1051), .B(KEYINPUT126), .C1(new_n827), .C2(new_n826), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1046), .A2(new_n1056), .A3(new_n832), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n1026), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1029), .B1(new_n1041), .B2(new_n1058), .ZN(G72));
  NAND2_X1  g873(.A1(new_n277), .A2(new_n287), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1036), .A2(new_n1021), .A3(new_n1039), .ZN(new_n1061));
  NAND2_X1  g875(.A1(G472), .A2(G902), .ZN(new_n1062));
  XOR2_X1   g876(.A(new_n1062), .B(KEYINPUT63), .Z(new_n1063));
  AOI21_X1  g877(.A(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n1046), .A2(new_n1056), .A3(new_n832), .A4(new_n1021), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n724), .B1(new_n1065), .B2(new_n1063), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n273), .A2(new_n301), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n925), .A2(new_n931), .A3(new_n1063), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1068), .A2(new_n977), .ZN(new_n1069));
  NOR3_X1   g883(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(G57));
endmodule


