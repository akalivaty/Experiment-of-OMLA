//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT81), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(G214), .B1(G237), .B2(G902), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(G210), .B1(G237), .B2(G902), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT82), .A2(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(G107), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(G101), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT85), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT82), .A2(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT82), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n203), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n198), .A2(KEYINPUT3), .A3(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n209), .B2(KEYINPUT3), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(G107), .A3(new_n200), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT83), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(new_n208), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G107), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n206), .B(new_n216), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT5), .A3(G119), .ZN(new_n226));
  INV_X1    g040(.A(G113), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT2), .B(G113), .Z(new_n229));
  AOI22_X1  g043(.A1(new_n224), .A2(new_n228), .B1(new_n229), .B2(new_n223), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n214), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n217), .B(KEYINPUT83), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n206), .B1(new_n233), .B2(new_n216), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G101), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n229), .B(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n231), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(new_n231), .C1(new_n235), .C2(new_n240), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(KEYINPUT6), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  INV_X1    g062(.A(G125), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n258), .A3(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT0), .A4(G128), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n249), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n255), .A2(KEYINPUT65), .A3(new_n258), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT65), .B1(new_n255), .B2(new_n258), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT91), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n252), .A2(new_n254), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT67), .B(G128), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(G143), .B2(new_n251), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n252), .A2(new_n254), .A3(new_n275), .A4(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G125), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n267), .A2(new_n272), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT92), .B(G224), .Z(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n284), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n267), .A2(new_n272), .A3(new_n286), .A4(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n246), .A2(new_n248), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n242), .B(KEYINPUT8), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n214), .A2(new_n222), .A3(new_n230), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n230), .B1(new_n214), .B2(new_n222), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT93), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(KEYINPUT93), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n267), .A2(new_n272), .A3(new_n281), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n265), .A2(new_n280), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n245), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n190), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n196), .B1(new_n290), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n300), .A2(new_n302), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n190), .A3(new_n195), .A4(new_n289), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n194), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G128), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n273), .B1(new_n276), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n278), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n214), .A2(new_n222), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT72), .B1(new_n277), .B2(new_n278), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT10), .A3(new_n222), .A4(new_n214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G134), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n324), .A3(new_n329), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n331), .B(KEYINPUT86), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n335), .B(new_n264), .C1(new_n268), .C2(new_n269), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(new_n238), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n236), .A2(G101), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT84), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n238), .A3(new_n336), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n235), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n319), .B(new_n333), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n335), .B1(new_n263), .B2(new_n264), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT84), .A3(new_n339), .A4(new_n238), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n341), .B2(new_n235), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n318), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n331), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI211_X1 g166(.A(KEYINPUT89), .B(new_n318), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n344), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G140), .ZN(new_n355));
  INV_X1    g169(.A(G953), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(G227), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n355), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT90), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n332), .B(new_n318), .C1(new_n348), .C2(new_n349), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n358), .ZN(new_n362));
  INV_X1    g176(.A(new_n358), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n344), .A2(KEYINPUT90), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n214), .A2(new_n222), .A3(new_n310), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n279), .B1(new_n214), .B2(new_n222), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT12), .B(new_n331), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n331), .B1(new_n365), .B2(new_n366), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n211), .A2(new_n212), .ZN(new_n373));
  AOI211_X1 g187(.A(KEYINPUT85), .B(new_n206), .C1(new_n209), .C2(new_n210), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n222), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n279), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n311), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(KEYINPUT87), .A3(KEYINPUT12), .A4(new_n331), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n369), .A2(new_n372), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n362), .A2(new_n364), .A3(new_n380), .ZN(new_n381));
  AOI211_X1 g195(.A(G469), .B(G902), .C1(new_n359), .C2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n344), .A2(new_n380), .A3(KEYINPUT88), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT88), .B1(new_n344), .B2(new_n380), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n358), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n344), .B(new_n363), .C1(new_n352), .C2(new_n353), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G469), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(G469), .A2(G902), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n192), .B(new_n307), .C1(new_n382), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n274), .A2(G119), .ZN(new_n392));
  INV_X1    g206(.A(G119), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT77), .B1(new_n393), .B2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT24), .B(G110), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(G128), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n393), .B2(G128), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT78), .B1(new_n399), .B2(KEYINPUT23), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n401), .A2(new_n402), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(G110), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n249), .A2(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT16), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n249), .A2(KEYINPUT16), .A3(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G146), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n408), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n405), .B(new_n411), .C1(G146), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n404), .A2(G110), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n409), .B2(new_n410), .ZN(new_n415));
  INV_X1    g229(.A(new_n411), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n392), .A2(new_n397), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n392), .B2(new_n394), .ZN(new_n418));
  OAI221_X1 g232(.A(new_n414), .B1(new_n415), .B2(new_n416), .C1(new_n418), .C2(new_n396), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G137), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n356), .A2(G221), .A3(G234), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n419), .A3(new_n423), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT80), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(G234), .B2(new_n190), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G902), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n425), .A2(new_n190), .A3(new_n426), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G472), .A2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n334), .A2(new_n336), .A3(new_n331), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT70), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n334), .A2(new_n447), .A3(new_n336), .A4(new_n331), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n321), .A2(new_n326), .A3(KEYINPUT66), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(G131), .C1(KEYINPUT66), .C2(new_n321), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n330), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(KEYINPUT71), .A3(new_n330), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n456), .B2(new_n316), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n239), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT68), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n376), .B2(new_n452), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n279), .A2(KEYINPUT68), .A3(new_n330), .A4(new_n451), .ZN(new_n462));
  INV_X1    g276(.A(new_n331), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n462), .C1(new_n270), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n459), .B1(new_n464), .B2(new_n449), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n239), .B1(new_n456), .B2(new_n316), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n446), .A2(new_n448), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT26), .B(G101), .Z(new_n469));
  NOR2_X1   g283(.A1(G237), .A2(G953), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G210), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT31), .B1(new_n466), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n474), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT75), .B(KEYINPUT28), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n464), .A2(new_n239), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT28), .B1(new_n467), .B2(new_n445), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n458), .A2(new_n465), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT31), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n468), .A4(new_n474), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT74), .ZN(new_n487));
  INV_X1    g301(.A(new_n475), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n485), .A4(new_n484), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n444), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n440), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n494), .B2(new_n442), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n446), .A2(new_n448), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n497), .A2(new_n467), .B1(new_n458), .B2(new_n465), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(new_n474), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n480), .A2(new_n477), .A3(new_n481), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT76), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n456), .A2(new_n316), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n446), .A2(new_n448), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n239), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n468), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n481), .B1(new_n505), .B2(KEYINPUT28), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n477), .A2(new_n496), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n484), .A2(new_n468), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n509), .B2(new_n477), .ZN(new_n510));
  INV_X1    g324(.A(new_n481), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n468), .A2(new_n479), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n474), .B(new_n511), .C1(new_n512), .C2(new_n478), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT76), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G472), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n439), .B1(new_n495), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n308), .A2(KEYINPUT67), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G128), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n521), .A3(G143), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n308), .A2(G143), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G134), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n325), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n225), .A2(G122), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n202), .B1(new_n529), .B2(KEYINPUT14), .ZN(new_n530));
  XNOR2_X1  g344(.A(G116), .B(G122), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n532), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n522), .B1(KEYINPUT13), .B2(new_n523), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n536), .A2(KEYINPUT97), .B1(KEYINPUT13), .B2(new_n523), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n522), .B(new_n538), .C1(KEYINPUT13), .C2(new_n523), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n325), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n531), .B(new_n202), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n527), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n189), .A2(G217), .A3(new_n356), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(new_n535), .C1(new_n540), .C2(new_n542), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n548), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n416), .B2(new_n415), .ZN(new_n554));
  INV_X1    g368(.A(new_n415), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT95), .A3(new_n411), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n470), .A2(G143), .A3(G214), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G143), .B1(new_n470), .B2(G214), .ZN(new_n559));
  OAI21_X1  g373(.A(G131), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n470), .A2(G214), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n253), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n329), .A3(new_n557), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n329), .B1(new_n562), .B2(new_n557), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n554), .A2(new_n556), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G113), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n198), .ZN(new_n570));
  XNOR2_X1  g384(.A(G125), .B(G140), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n251), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT18), .B(G131), .C1(new_n558), .C2(new_n559), .ZN(new_n573));
  NAND2_X1  g387(.A1(KEYINPUT18), .A2(G131), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n562), .A2(new_n557), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n568), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n568), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n190), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT96), .B(G475), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT20), .ZN(new_n582));
  INV_X1    g396(.A(new_n570), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n558), .A2(new_n559), .A3(G131), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n411), .B1(new_n584), .B2(new_n566), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT19), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n412), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n571), .A2(KEYINPUT19), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n251), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n592), .A3(new_n251), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n585), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n576), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n568), .A2(new_n570), .A3(new_n576), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(G475), .A2(G902), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n599), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT20), .B(new_n601), .C1(new_n596), .C2(new_n597), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n581), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(G234), .A2(G237), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G952), .A3(new_n356), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(G902), .A3(G953), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT98), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT21), .B(G898), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n552), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n391), .A2(new_n518), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT99), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  AND2_X1   g429(.A1(new_n387), .A2(new_n388), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n359), .A2(new_n381), .ZN(new_n617));
  INV_X1    g431(.A(G469), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n190), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n191), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n493), .B2(new_n190), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n441), .B1(new_n483), .B2(new_n491), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n622), .A2(new_n623), .A3(new_n439), .ZN(new_n624));
  INV_X1    g438(.A(new_n611), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n307), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n545), .A2(new_n547), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n545), .A2(new_n629), .A3(new_n547), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(G478), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n549), .A2(new_n190), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n548), .B2(new_n549), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n603), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n620), .A2(new_n624), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NAND2_X1  g453(.A1(new_n493), .A2(new_n190), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  INV_X1    g455(.A(new_n439), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n494), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n192), .B1(new_n382), .B2(new_n389), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n551), .A2(new_n603), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n307), .A2(new_n625), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n307), .A2(KEYINPUT100), .A3(new_n625), .A4(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT101), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n424), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n420), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n431), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n438), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(new_n612), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n641), .A2(new_n494), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n390), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT37), .B(G110), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  INV_X1    g478(.A(new_n307), .ZN(new_n665));
  INV_X1    g479(.A(new_n646), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n493), .A2(new_n443), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(KEYINPUT32), .B2(new_n623), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n514), .B1(new_n510), .B2(new_n513), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n497), .A2(new_n467), .B1(new_n503), .B2(new_n239), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT28), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n511), .B(new_n507), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n190), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n621), .B1(new_n675), .B2(new_n515), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n667), .B(new_n659), .C1(new_n669), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n605), .B(KEYINPUT102), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(new_n609), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n192), .B(new_n682), .C1(new_n382), .C2(new_n389), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n308), .ZN(G30));
  XOR2_X1   g499(.A(new_n681), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n620), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n190), .B1(new_n505), .B2(new_n474), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n498), .A2(new_n477), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n668), .B(new_n692), .C1(KEYINPUT32), .C2(new_n623), .ZN(new_n693));
  INV_X1    g507(.A(new_n659), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n304), .A2(new_n306), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT38), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n552), .A2(new_n603), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n695), .A2(new_n697), .A3(new_n194), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n688), .A2(new_n689), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  NAND2_X1  g515(.A1(new_n494), .A2(new_n442), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n668), .A3(new_n517), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n603), .A2(new_n631), .A3(new_n633), .A4(new_n682), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n634), .A2(new_n706), .A3(new_n603), .A4(new_n682), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n665), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n620), .A2(new_n703), .A3(new_n659), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(new_n380), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n344), .A2(new_n363), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n360), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n364), .A2(new_n714), .B1(new_n354), .B2(new_n358), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n192), .A3(new_n619), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n518), .A2(new_n636), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n518), .A2(new_n651), .A3(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND4_X1  g536(.A1(new_n717), .A2(new_n307), .A3(new_n703), .A4(new_n660), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n192), .A3(new_n619), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n626), .A3(new_n698), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n483), .B2(new_n491), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(new_n621), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n476), .A2(new_n482), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n490), .B2(new_n487), .ZN(new_n732));
  OAI211_X1 g546(.A(KEYINPUT104), .B(G472), .C1(new_n732), .C2(G902), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n506), .A2(new_n474), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n485), .B1(new_n488), .B2(new_n484), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n490), .B2(new_n487), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n441), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n727), .A2(new_n734), .A3(new_n642), .A4(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n730), .B2(new_n733), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n727), .B1(new_n741), .B2(new_n642), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n726), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AND3_X1   g558(.A1(new_n705), .A2(new_n707), .A3(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT106), .B1(new_n705), .B2(new_n707), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n725), .A2(new_n747), .A3(new_n665), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n694), .B(new_n738), .C1(new_n730), .C2(new_n733), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  OAI21_X1  g565(.A(KEYINPUT107), .B1(new_n732), .B2(new_n444), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n492), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n702), .A2(new_n517), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n642), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n619), .A2(new_n388), .A3(new_n387), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n708), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n705), .A2(new_n707), .A3(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n191), .A2(new_n194), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n304), .A2(new_n306), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n757), .A2(new_n761), .A3(KEYINPUT42), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT108), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n764), .B1(new_n382), .B2(new_n389), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT42), .B1(new_n745), .B2(new_n746), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n642), .A4(new_n755), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n763), .B1(new_n616), .B2(new_n619), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n518), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n766), .A2(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n329), .ZN(G33));
  NOR2_X1   g590(.A1(new_n666), .A2(new_n681), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n518), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  NAND2_X1  g593(.A1(new_n385), .A2(new_n386), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n385), .A2(KEYINPUT45), .A3(new_n386), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n388), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT46), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n788));
  OAI221_X1 g602(.A(new_n619), .B1(KEYINPUT46), .B2(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n192), .ZN(new_n790));
  INV_X1    g604(.A(new_n634), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n603), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n603), .B2(KEYINPUT110), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n792), .B(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n659), .C1(new_n623), .C2(new_n622), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT44), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n696), .A2(new_n194), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT111), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n790), .A2(new_n686), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(new_n798), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n439), .A2(new_n707), .A3(new_n705), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n703), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  INV_X1    g624(.A(new_n626), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n646), .B(KEYINPUT113), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n620), .A2(new_n624), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n721), .A2(new_n723), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n703), .A2(new_n642), .A3(new_n612), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n391), .B1(new_n645), .B2(new_n636), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n642), .B1(new_n669), .B2(new_n676), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n725), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n662), .B1(new_n818), .B2(new_n636), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n814), .A2(new_n743), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n767), .A2(new_n747), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n749), .A2(new_n821), .A3(KEYINPUT114), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT104), .B1(new_n640), .B2(G472), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n729), .A2(new_n728), .A3(new_n621), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n659), .B(new_n739), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n757), .A2(new_n761), .A3(new_n764), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n552), .A2(new_n603), .A3(new_n681), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n798), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n620), .A2(new_n703), .A3(new_n659), .A4(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n778), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n820), .A2(new_n775), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n618), .B1(new_n617), .B2(new_n190), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n382), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n192), .A3(new_n761), .A4(new_n307), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n839), .A2(new_n826), .B1(new_n677), .B2(new_n683), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n659), .B1(new_n669), .B2(new_n676), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n644), .ZN(new_n843));
  INV_X1    g657(.A(new_n683), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n665), .A2(new_n698), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n693), .A2(new_n845), .A3(new_n694), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n843), .A2(new_n709), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n836), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n844), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n710), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(new_n840), .A3(KEYINPUT52), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n835), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n390), .A2(new_n661), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n613), .A2(new_n854), .A3(new_n718), .A4(new_n637), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n721), .A2(new_n723), .A3(new_n813), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n766), .A2(new_n771), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n774), .A2(new_n772), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n778), .A2(new_n832), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n828), .B2(new_n822), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n860), .A3(new_n862), .A4(new_n743), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n841), .A2(new_n847), .A3(new_n836), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT52), .B1(new_n850), .B2(new_n840), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n853), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT115), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n693), .A2(new_n439), .A3(new_n605), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n725), .A2(new_n803), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT117), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n880), .A2(new_n603), .A3(new_n634), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n795), .A2(new_n679), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n749), .A2(new_n882), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n742), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n741), .A2(new_n727), .A3(new_n642), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n882), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n717), .A2(new_n194), .A3(new_n697), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT50), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(KEYINPUT50), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(new_n838), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n192), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n807), .A2(new_n808), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n889), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n799), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n885), .B(new_n896), .C1(new_n899), .C2(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n900), .A2(new_n665), .A3(new_n725), .ZN(new_n904));
  INV_X1    g718(.A(new_n756), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n882), .A3(new_n878), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT48), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G952), .A3(new_n356), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n880), .A2(new_n635), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n904), .A2(new_n908), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n913));
  INV_X1    g727(.A(new_n898), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n806), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n884), .B1(new_n915), .B2(new_n901), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n895), .B(KEYINPUT116), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n903), .B(new_n912), .C1(new_n918), .C2(KEYINPUT51), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n876), .A2(new_n919), .B1(G952), .B2(G953), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n642), .A2(new_n762), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT112), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n697), .A3(new_n792), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n897), .A2(KEYINPUT49), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n693), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(KEYINPUT49), .B2(new_n897), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n926), .ZN(G75));
  OR2_X1    g741(.A1(new_n356), .A2(G952), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT119), .Z(new_n929));
  NOR2_X1   g743(.A1(new_n869), .A2(new_n190), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n930), .B2(G210), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n246), .A2(new_n248), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n288), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n929), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT118), .B1(new_n869), .B2(new_n190), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n196), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n939), .B2(new_n941), .ZN(G51));
  INV_X1    g756(.A(new_n929), .ZN(new_n943));
  INV_X1    g757(.A(new_n784), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n937), .A2(new_n944), .A3(new_n938), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT120), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n388), .B(KEYINPUT57), .Z(new_n947));
  NAND3_X1  g761(.A1(new_n870), .A2(new_n871), .A3(new_n947), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n945), .A2(KEYINPUT120), .B1(new_n948), .B2(new_n617), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n946), .B2(new_n949), .ZN(G54));
  NAND2_X1  g764(.A1(new_n937), .A2(new_n938), .ZN(new_n951));
  NAND2_X1  g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n951), .A2(new_n598), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n598), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(G60));
  NAND2_X1  g769(.A1(new_n628), .A2(new_n630), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT121), .Z(new_n957));
  XOR2_X1   g771(.A(new_n632), .B(KEYINPUT59), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n929), .B1(new_n872), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(KEYINPUT122), .B(new_n929), .C1(new_n872), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n957), .B1(new_n876), .B2(new_n958), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G63));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n853), .B2(new_n868), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n864), .B1(new_n863), .B2(new_n867), .ZN(new_n974));
  INV_X1    g788(.A(new_n820), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n834), .A2(new_n775), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n970), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n657), .B(KEYINPUT124), .Z(new_n981));
  AOI21_X1  g795(.A(KEYINPUT125), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT123), .B1(new_n978), .B2(new_n970), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n972), .B(new_n969), .C1(new_n974), .C2(new_n977), .ZN(new_n984));
  OAI211_X1 g798(.A(KEYINPUT125), .B(new_n981), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n967), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n983), .A2(new_n984), .ZN(new_n988));
  INV_X1    g802(.A(new_n428), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n943), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n982), .B2(new_n986), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI221_X1 g807(.A(new_n990), .B1(new_n967), .B2(KEYINPUT61), .C1(new_n982), .C2(new_n986), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n283), .B2(new_n610), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n975), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n932), .B1(G898), .B2(new_n356), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT127), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(G69));
  INV_X1    g814(.A(new_n809), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n790), .A2(new_n686), .A3(new_n905), .A4(new_n845), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n840), .B1(new_n843), .B2(new_n709), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n860), .A2(new_n1003), .A3(new_n778), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n801), .A3(new_n1004), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n1001), .A2(G953), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n464), .A2(new_n449), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n458), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n589), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(G900), .B2(G953), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n812), .B1(new_n603), .B2(new_n634), .ZN(new_n1011));
  OR4_X1    g825(.A1(new_n817), .A2(new_n687), .A3(new_n803), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1003), .A2(new_n700), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT62), .Z(new_n1014));
  NAND4_X1  g828(.A1(new_n809), .A2(new_n801), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n356), .ZN(new_n1016));
  AOI22_X1  g830(.A1(new_n1006), .A2(new_n1010), .B1(new_n1016), .B2(new_n1009), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n356), .B1(G227), .B2(G900), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1017), .B(new_n1019), .ZN(G72));
  NOR2_X1   g834(.A1(new_n1015), .A2(new_n820), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT63), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n691), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1001), .A2(new_n1005), .A3(new_n820), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n477), .B(new_n498), .C1(new_n1025), .C2(new_n1023), .ZN(new_n1026));
  AOI22_X1  g840(.A1(new_n509), .A2(new_n477), .B1(new_n488), .B2(new_n484), .ZN(new_n1027));
  OR3_X1    g841(.A1(new_n869), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n929), .A2(new_n1024), .A3(new_n1026), .A4(new_n1028), .ZN(G57));
endmodule


