//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1155, new_n1156, new_n1158, new_n1159,
    new_n1160, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222, new_n1223;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT65), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n252), .B(KEYINPUT67), .Z(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G226), .ZN(new_n254));
  INV_X1    g0054(.A(new_n251), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(new_n250), .A3(G274), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n258), .A2(new_n259), .B1(new_n225), .B2(new_n257), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n260), .B1(G222), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n254), .B(new_n256), .C1(new_n267), .C2(new_n250), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT71), .B(G200), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n215), .B1(new_n209), .B2(new_n261), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(new_n207), .A3(G1), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n206), .A2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G50), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n275), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(G50), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n273), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n207), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(G150), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n268), .A2(new_n294), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n272), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n268), .A2(G179), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT68), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n289), .B1(new_n268), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n257), .A2(G232), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n307), .B1(new_n227), .B2(new_n257), .C1(new_n258), .C2(new_n220), .ZN(new_n308));
  INV_X1    g0108(.A(new_n250), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n253), .A2(G244), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n256), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  INV_X1    g0116(.A(new_n285), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n282), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n319), .B1(new_n207), .B2(new_n225), .C1(new_n283), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n273), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n276), .A2(G77), .A3(new_n277), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(G77), .C2(new_n279), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n312), .A2(new_n301), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n315), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n312), .B2(new_n269), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G190), .B2(new_n313), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n312), .A2(new_n328), .A3(new_n294), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n330), .A2(new_n331), .A3(new_n324), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n304), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n282), .B1(new_n206), .B2(G20), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n276), .A2(new_n334), .B1(new_n275), .B2(new_n282), .ZN(new_n335));
  INV_X1    g0135(.A(G58), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n219), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n337), .B2(new_n201), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n285), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n265), .B2(new_n207), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n342), .B(G20), .C1(new_n262), .C2(new_n264), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT77), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n342), .B1(new_n257), .B2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n219), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT77), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT16), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n340), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n273), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n335), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n306), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n309), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n256), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n361), .A2(new_n363), .A3(new_n314), .ZN(new_n364));
  AOI21_X1  g0164(.A(G169), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n301), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(new_n363), .A3(new_n314), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n355), .A2(new_n356), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n356), .B1(new_n355), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT79), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G190), .B2(new_n367), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n335), .C1(new_n351), .C2(new_n354), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT80), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n335), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n352), .B1(new_n349), .B2(KEYINPUT77), .ZN(new_n388));
  AOI211_X1 g0188(.A(new_n345), .B(new_n219), .C1(new_n347), .C2(new_n348), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n349), .A2(new_n340), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n281), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n385), .B1(new_n393), .B2(new_n378), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT81), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n379), .B1(new_n384), .B2(new_n382), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n393), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT81), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n366), .A2(new_n371), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n400), .B2(new_n393), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT79), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n355), .A2(new_n356), .A3(new_n372), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n375), .A2(new_n395), .A3(new_n399), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n266), .A2(G226), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT74), .ZN(new_n408));
  INV_X1    g0208(.A(G97), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n261), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n305), .B2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n309), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n253), .A2(G238), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n256), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n250), .B1(new_n408), .B2(new_n411), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT13), .B1(new_n419), .B2(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G179), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n413), .B2(new_n417), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n419), .A2(KEYINPUT13), .A3(new_n416), .ZN(new_n423));
  OAI21_X1  g0223(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(KEYINPUT14), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT14), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n301), .B1(new_n418), .B2(new_n420), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT75), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n425), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n276), .A2(G68), .A3(new_n277), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n275), .A2(new_n219), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT11), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n225), .B2(new_n283), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n273), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n432), .B(new_n434), .C1(new_n435), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n435), .B2(new_n438), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT76), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n422), .A2(new_n423), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G190), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n440), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n376), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n333), .A2(new_n406), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n257), .A2(G257), .A3(new_n306), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n452), .B1(new_n453), .B2(new_n257), .C1(new_n258), .C2(new_n228), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT89), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n309), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n250), .A2(G274), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT5), .B(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n309), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G270), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n207), .C1(G33), .C2(new_n409), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n273), .B(new_n467), .C1(new_n207), .C2(G116), .ZN(new_n468));
  XOR2_X1   g0268(.A(new_n468), .B(KEYINPUT20), .Z(new_n469));
  NOR2_X1   g0269(.A1(new_n279), .A2(G116), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n276), .B1(G1), .B2(new_n261), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(G116), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n301), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT21), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n465), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n469), .A2(new_n473), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n465), .B2(G200), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n294), .B2(new_n465), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n464), .A2(G179), .A3(new_n462), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n480), .A2(new_n457), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT6), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(KEYINPUT6), .B2(new_n409), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT82), .B(G107), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n491), .A2(KEYINPUT83), .ZN(new_n492));
  OAI21_X1  g0292(.A(G107), .B1(new_n341), .B2(new_n343), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(KEYINPUT83), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n273), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n471), .A2(G97), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G97), .B2(new_n275), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n497), .B(KEYINPUT84), .C1(G97), .C2(new_n275), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n466), .C1(new_n222), .C2(new_n258), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT4), .B1(new_n266), .B2(G244), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n309), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n463), .A2(G257), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n462), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n301), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G179), .B2(new_n509), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n495), .A2(new_n273), .B1(new_n500), .B2(new_n501), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(G200), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n507), .A2(new_n508), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(G190), .A3(new_n462), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n257), .A2(new_n207), .A3(G87), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n261), .A2(new_n521), .A3(G20), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n207), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n227), .A2(KEYINPUT23), .A3(G20), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT24), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n273), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT25), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n279), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n227), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n472), .A2(G107), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n257), .A2(new_n306), .ZN(new_n537));
  OAI221_X1 g0337(.A(new_n535), .B1(new_n261), .B2(new_n536), .C1(new_n537), .C2(new_n222), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n309), .B1(G264), .B2(new_n463), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n462), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G179), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n301), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n513), .A2(new_n518), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n257), .A2(new_n207), .A3(G68), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n283), .A2(new_n409), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(KEYINPUT19), .B2(new_n547), .ZN(new_n548));
  XOR2_X1   g0348(.A(KEYINPUT86), .B(G87), .Z(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n486), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT87), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(new_n410), .B2(KEYINPUT19), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n548), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n320), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n554), .A2(new_n281), .B1(new_n279), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(G87), .B2(new_n472), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n458), .A2(new_n460), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n250), .B(G250), .C1(G1), .C2(new_n459), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n258), .A2(new_n226), .B1(new_n261), .B2(new_n521), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n266), .A2(new_n561), .A3(G238), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT85), .B1(new_n537), .B2(new_n220), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n558), .B(new_n559), .C1(new_n564), .C2(new_n250), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT88), .ZN(new_n568));
  OR3_X1    g0368(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n294), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n565), .A2(new_n269), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n557), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n301), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n471), .A2(new_n320), .ZN(new_n573));
  OAI221_X1 g0373(.A(new_n572), .B1(G179), .B2(new_n565), .C1(new_n556), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n540), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n540), .A2(G200), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR3_X1    g0379(.A1(new_n534), .A2(KEYINPUT90), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT90), .B1(new_n534), .B2(new_n579), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND4_X1   g0382(.A1(new_n451), .A2(new_n485), .A3(new_n545), .A4(new_n582), .ZN(G372));
  NOR2_X1   g0383(.A1(new_n373), .A2(new_n374), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n446), .A2(new_n447), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n443), .B1(new_n585), .B2(new_n327), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n395), .A2(new_n399), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n513), .A2(new_n518), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n580), .A2(new_n581), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n479), .A2(new_n484), .A3(new_n543), .ZN(new_n592));
  INV_X1    g0392(.A(new_n556), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n472), .A2(G87), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n567), .A3(new_n570), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n574), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT26), .B1(new_n575), .B2(new_n513), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n514), .A2(new_n511), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n574), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n589), .B1(new_n450), .B2(new_n604), .ZN(G369));
  NAND3_X1  g0405(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n606), .A2(KEYINPUT27), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(KEYINPUT27), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(G213), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g0409(.A(new_n609), .B(KEYINPUT91), .Z(new_n610));
  INV_X1    g0410(.A(KEYINPUT92), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n611), .A2(G343), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(G343), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n480), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n485), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n479), .A2(new_n484), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G330), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n534), .A2(new_n616), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT93), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n591), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n543), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n534), .A2(new_n542), .A3(new_n615), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n625), .A2(new_n626), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n619), .A2(new_n616), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n626), .A3(new_n632), .ZN(G399));
  NOR2_X1   g0433(.A1(new_n551), .A2(G116), .ZN(new_n634));
  INV_X1    g0434(.A(new_n210), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G41), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(G1), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT94), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n213), .B2(new_n637), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT28), .Z(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT26), .B1(new_n513), .B2(new_n596), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n574), .B(KEYINPUT96), .Z(new_n644));
  NAND4_X1  g0444(.A1(new_n600), .A2(new_n601), .A3(new_n574), .A4(new_n571), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n597), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n616), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT29), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n604), .A2(new_n616), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n516), .A2(new_n483), .A3(new_n539), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n457), .A2(new_n566), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT30), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n566), .A2(new_n576), .A3(G179), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n465), .A3(new_n509), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n660), .A2(KEYINPUT31), .A3(new_n616), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT31), .B1(new_n660), .B2(new_n616), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n582), .A2(new_n545), .A3(new_n485), .A4(new_n615), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n642), .B1(new_n668), .B2(G1), .ZN(G364));
  NOR2_X1   g0469(.A1(new_n274), .A2(G20), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n206), .B1(new_n670), .B2(G45), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n636), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n635), .A2(new_n257), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n214), .B2(new_n459), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n459), .B2(new_n247), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n635), .A2(new_n265), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(G355), .B1(new_n521), .B2(new_n635), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(G13), .A2(G33), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT97), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n207), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT98), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n215), .B1(G20), .B2(new_n301), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n674), .B1(new_n681), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  NOR2_X1   g0491(.A1(new_n207), .A2(new_n314), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G200), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G190), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(KEYINPUT33), .B(G317), .Z(new_n696));
  NOR2_X1   g0496(.A1(new_n693), .A2(new_n294), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G326), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G190), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n207), .A2(G179), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n701), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(G311), .A2(new_n703), .B1(new_n706), .B2(G329), .ZN(new_n707));
  INV_X1    g0507(.A(G322), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n376), .A2(G190), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n709), .A2(new_n207), .A3(new_n314), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n707), .B(new_n265), .C1(new_n708), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n269), .A2(G190), .A3(new_n704), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n700), .B(new_n712), .C1(G303), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G283), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n269), .A2(new_n294), .A3(new_n704), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT100), .Z(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(G20), .B1(new_n709), .B2(G179), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT101), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI221_X1 g0524(.A(new_n715), .B1(new_n716), .B2(new_n719), .C1(new_n536), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G50), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n698), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n706), .A2(G159), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n695), .A2(new_n219), .B1(new_n728), .B2(KEYINPUT32), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n727), .B(new_n729), .C1(KEYINPUT32), .C2(new_n728), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n718), .A2(G107), .ZN(new_n731));
  INV_X1    g0531(.A(new_n724), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G97), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n257), .B1(new_n702), .B2(new_n225), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n713), .A2(new_n549), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n734), .B(new_n735), .C1(G58), .C2(new_n710), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n730), .A2(new_n731), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n725), .A2(KEYINPUT102), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT102), .B1(new_n725), .B2(new_n737), .ZN(new_n739));
  INV_X1    g0539(.A(new_n688), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n691), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n620), .B2(new_n686), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n621), .A2(new_n674), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n620), .A2(G330), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT103), .ZN(G396));
  AND2_X1   g0547(.A1(new_n324), .A2(new_n616), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n326), .B1(new_n332), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n327), .A2(new_n615), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n650), .B(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n673), .B1(new_n752), .B2(new_n667), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n667), .B2(new_n752), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n716), .A2(new_n695), .B1(new_n698), .B2(new_n453), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n265), .B1(new_n711), .B2(new_n536), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n702), .A2(new_n521), .B1(new_n705), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n718), .A2(G87), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n714), .A2(G107), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n759), .A2(new_n733), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G132), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n257), .B1(new_n705), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n714), .B2(G50), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n703), .A2(G159), .B1(new_n710), .B2(G143), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  INV_X1    g0567(.A(G150), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n766), .B1(new_n698), .B2(new_n767), .C1(new_n768), .C2(new_n695), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT34), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n765), .B1(new_n336), .B2(new_n724), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n718), .A2(G68), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n762), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n688), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n688), .A2(new_n682), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n674), .B1(new_n225), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n778), .C1(new_n751), .C2(new_n683), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n754), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G384));
  INV_X1    g0581(.A(new_n490), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT35), .ZN(new_n783));
  OAI211_X1 g0583(.A(G116), .B(new_n216), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT36), .ZN(new_n786));
  OR3_X1    g0586(.A1(new_n213), .A2(new_n225), .A3(new_n337), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n726), .A2(G68), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n206), .B(G13), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n335), .B1(new_n354), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n610), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n405), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT105), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n372), .A2(new_n792), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n379), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT37), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT104), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n355), .A2(new_n372), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n355), .A2(new_n610), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT37), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n379), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT104), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n798), .A2(new_n805), .A3(KEYINPUT37), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n800), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT38), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n804), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n405), .A2(new_n794), .B1(new_n809), .B2(new_n800), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n808), .B1(KEYINPUT38), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n796), .B1(new_n810), .B2(KEYINPUT38), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT39), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT39), .ZN(new_n814));
  INV_X1    g0614(.A(new_n610), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n393), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n401), .B(new_n403), .C1(new_n383), .C2(new_n394), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n379), .B1(new_n400), .B2(new_n393), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT37), .B1(new_n818), .B2(new_n816), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n804), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT107), .B1(new_n820), .B2(KEYINPUT38), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(KEYINPUT38), .B2(new_n810), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT107), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n823), .A2(new_n795), .A3(KEYINPUT38), .A4(new_n807), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT108), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n813), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n813), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n431), .A2(new_n442), .A3(new_n616), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n584), .A2(new_n610), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT106), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n811), .B2(new_n812), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n795), .A2(new_n807), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT105), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT106), .A4(new_n808), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n441), .A2(new_n616), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n585), .B(new_n841), .C1(new_n431), .C2(new_n442), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n427), .A2(new_n430), .ZN(new_n843));
  INV_X1    g0643(.A(new_n425), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n441), .B(new_n616), .C1(new_n845), .C2(new_n448), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n751), .B(new_n615), .C1(new_n598), .C2(new_n603), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n750), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n832), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n831), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n589), .B1(new_n450), .B2(new_n652), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n842), .A2(new_n846), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n665), .A3(new_n751), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n834), .B2(new_n839), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT40), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n854), .A2(new_n751), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n822), .A2(new_n824), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT40), .A4(new_n665), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n451), .A2(new_n665), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(G330), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n206), .B2(new_n670), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n853), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n790), .B1(new_n867), .B2(new_n868), .ZN(G367));
  OAI21_X1  g0669(.A(new_n590), .B1(new_n514), .B2(new_n615), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n870), .A2(new_n543), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n616), .B1(new_n871), .B2(new_n513), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT42), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n870), .B1(new_n513), .B2(new_n615), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n632), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n630), .A2(KEYINPUT42), .A3(new_n631), .A4(new_n874), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n557), .A2(new_n615), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT109), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n597), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n574), .B2(new_n880), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT110), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT43), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(KEYINPUT43), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n878), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n628), .A2(new_n874), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n890), .B(new_n891), .Z(new_n892));
  XOR2_X1   g0692(.A(new_n636), .B(KEYINPUT41), .Z(new_n893));
  AOI21_X1  g0693(.A(new_n874), .B1(new_n632), .B2(new_n626), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(KEYINPUT44), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(KEYINPUT44), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n632), .A2(new_n626), .A3(new_n874), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT45), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n900), .A3(new_n629), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n895), .A2(new_n896), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n628), .B1(new_n902), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n627), .B1(new_n619), .B2(new_n616), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n632), .A2(new_n621), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n621), .B1(new_n632), .B2(new_n904), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n668), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT111), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n908), .A2(KEYINPUT111), .A3(new_n668), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n901), .A2(new_n903), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n893), .B1(new_n913), .B2(new_n668), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n892), .B1(new_n914), .B2(new_n672), .ZN(new_n915));
  INV_X1    g0715(.A(new_n689), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n676), .A2(new_n239), .B1(new_n210), .B2(new_n320), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n673), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n703), .A2(G50), .B1(new_n710), .B2(G150), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n257), .C1(new_n767), .C2(new_n705), .ZN(new_n920));
  INV_X1    g0720(.A(G143), .ZN(new_n921));
  INV_X1    g0721(.A(G159), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n921), .A2(new_n698), .B1(new_n695), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n924), .B1(new_n336), .B2(new_n713), .C1(new_n225), .C2(new_n717), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n724), .A2(new_n219), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G294), .A2(new_n694), .B1(new_n697), .B2(G311), .ZN(new_n927));
  INV_X1    g0727(.A(new_n717), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(G97), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n257), .B1(new_n706), .B2(G317), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n703), .A2(G283), .B1(new_n710), .B2(G303), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n927), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n714), .A2(KEYINPUT46), .A3(G116), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT46), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n713), .B2(new_n521), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(new_n724), .C2(new_n227), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n925), .A2(new_n926), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT47), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n918), .B1(new_n938), .B2(new_n688), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n882), .B2(new_n686), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n915), .A2(new_n940), .ZN(G387));
  OAI21_X1  g0741(.A(new_n636), .B1(new_n908), .B2(new_n668), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n911), .B2(new_n912), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n265), .B1(new_n705), .B2(new_n699), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n703), .A2(G303), .B1(new_n710), .B2(G317), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n698), .B2(new_n708), .C1(new_n757), .C2(new_n695), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT48), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n716), .B2(new_n724), .C1(new_n536), .C2(new_n713), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT49), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n944), .B(new_n952), .C1(G116), .C2(new_n928), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n711), .A2(new_n726), .B1(new_n705), .B2(new_n768), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n265), .B(new_n954), .C1(G68), .C2(new_n703), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n732), .A2(new_n555), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n714), .A2(G77), .ZN(new_n957));
  INV_X1    g0757(.A(new_n282), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G159), .A2(new_n697), .B1(new_n694), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G97), .B2(new_n718), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n688), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n634), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n679), .B1(new_n227), .B2(new_n635), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n958), .A2(KEYINPUT50), .A3(new_n726), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT50), .B1(new_n958), .B2(new_n726), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n459), .B1(new_n219), .B2(new_n225), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n675), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n236), .A2(new_n459), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n916), .B1(new_n970), .B2(KEYINPUT112), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT112), .B2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n962), .A2(new_n673), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n627), .B2(new_n687), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n908), .B2(new_n672), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n943), .A2(new_n976), .ZN(G393));
  INV_X1    g0777(.A(new_n903), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n902), .A2(new_n899), .A3(new_n628), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n978), .A2(new_n979), .A3(new_n671), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n875), .A2(new_n687), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n689), .B1(new_n409), .B2(new_n210), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n244), .A2(new_n675), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n673), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n697), .A2(G317), .B1(G311), .B2(new_n710), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT52), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT113), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n713), .A2(new_n716), .B1(new_n708), .B2(new_n705), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n257), .B1(new_n703), .B2(G294), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n988), .A2(new_n987), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n731), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n724), .A2(new_n521), .B1(new_n453), .B2(new_n695), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT114), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n698), .A2(new_n768), .B1(new_n922), .B2(new_n711), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT51), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G77), .B2(new_n732), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n996), .B2(new_n995), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n713), .A2(new_n219), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n257), .B1(new_n705), .B2(new_n921), .C1(new_n282), .C2(new_n702), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G50), .C2(new_n694), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n760), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n992), .A2(new_n994), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n984), .B1(new_n1004), .B2(new_n688), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n980), .B1(new_n981), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n911), .A2(new_n912), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n979), .B2(new_n978), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n636), .A3(new_n913), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(G390));
  NAND4_X1  g0810(.A1(new_n666), .A2(new_n406), .A3(new_n449), .A4(new_n333), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n589), .B(new_n1011), .C1(new_n652), .C2(new_n450), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n848), .A2(new_n750), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n858), .A2(new_n666), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n854), .B1(new_n666), .B2(new_n751), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n648), .A2(new_n749), .B1(new_n327), .B2(new_n615), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n666), .A2(new_n751), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1014), .C1(new_n1019), .C2(new_n854), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1012), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1013), .A2(new_n854), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n830), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n827), .B2(new_n828), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n859), .C1(new_n1018), .C2(new_n847), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1014), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1014), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1022), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n849), .A2(new_n830), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n813), .A2(new_n825), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT108), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n813), .A2(new_n825), .A3(new_n826), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1027), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1015), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n1030), .A3(new_n1021), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1032), .A2(new_n636), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT117), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1027), .A2(new_n1014), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n672), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1045), .B2(new_n1028), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n671), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1039), .A2(new_n1047), .A3(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n711), .A2(new_n521), .B1(new_n702), .B2(new_n409), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n227), .A2(new_n695), .B1(new_n698), .B2(new_n716), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(G294), .C2(new_n706), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n773), .C1(new_n225), .C2(new_n724), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n265), .B1(new_n713), .B2(new_n221), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT54), .B(G143), .ZN(new_n1056));
  INV_X1    g0856(.A(G125), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n702), .A2(new_n1056), .B1(new_n705), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n265), .B(new_n1058), .C1(G132), .C2(new_n710), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G128), .A2(new_n697), .B1(new_n694), .B2(G137), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n726), .B2(new_n717), .C1(new_n922), .C2(new_n724), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n714), .A2(G150), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT53), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1053), .A2(new_n1055), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n688), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n674), .B1(new_n282), .B2(new_n777), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n829), .C2(new_n683), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1042), .B1(new_n1049), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1068), .ZN(new_n1070));
  AOI211_X1 g0870(.A(KEYINPUT117), .B(new_n1070), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1041), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT118), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(KEYINPUT118), .B(new_n1041), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(G378));
  NOR2_X1   g0877(.A1(new_n289), .A2(new_n815), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n304), .B(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1079), .B(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n857), .A2(G330), .A3(new_n860), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1082), .ZN(new_n1084));
  OAI211_X1 g0884(.A(G330), .B(new_n860), .C1(new_n856), .C2(KEYINPUT40), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n1086), .A3(new_n831), .A4(new_n850), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n851), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1012), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1087), .A2(new_n1090), .B1(new_n1040), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT120), .B1(new_n1092), .B2(KEYINPUT57), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n637), .B1(new_n1092), .B2(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1090), .A2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1040), .A2(new_n1091), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT120), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT57), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1093), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1084), .A2(new_n684), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n409), .A2(new_n695), .B1(new_n698), .B2(new_n521), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n711), .A2(new_n227), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n257), .A2(G41), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n702), .A2(new_n320), .B1(new_n705), .B2(new_n716), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n926), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n928), .A2(G58), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n957), .A4(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT58), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1105), .B(new_n726), .C1(G33), .C2(G41), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n703), .A2(G137), .B1(new_n710), .B2(G128), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1057), .B2(new_n698), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G132), .B2(new_n694), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n768), .B2(new_n724), .C1(new_n713), .C2(new_n1056), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n928), .A2(G159), .ZN(new_n1118));
  AOI211_X1 g0918(.A(G33), .B(G41), .C1(new_n706), .C2(G124), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1111), .B(new_n1112), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT119), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n740), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n674), .B(new_n1126), .C1(new_n726), .C2(new_n777), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1095), .A2(new_n672), .B1(new_n1102), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1101), .A2(new_n1128), .ZN(G375));
  NAND2_X1  g0929(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1012), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n893), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1022), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n847), .A2(new_n682), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT121), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n724), .A2(new_n726), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1109), .B1(new_n922), .B2(new_n713), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n763), .A2(new_n698), .B1(new_n695), .B2(new_n1056), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n706), .A2(G128), .B1(new_n710), .B2(G137), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n257), .C1(new_n768), .C2(new_n702), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n702), .A2(new_n227), .B1(new_n705), .B2(new_n453), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n257), .B(new_n1143), .C1(G283), .C2(new_n710), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n714), .A2(G97), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G116), .A2(new_n694), .B1(new_n697), .B2(G294), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(new_n956), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G77), .B2(new_n718), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n688), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n674), .B1(new_n219), .B2(new_n777), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1136), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1131), .B2(new_n671), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1134), .A2(new_n1153), .ZN(G381));
  OR3_X1    g0954(.A1(new_n943), .A2(G396), .A3(new_n976), .ZN(new_n1155));
  OR4_X1    g0955(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1155), .ZN(new_n1156));
  OR4_X1    g0956(.A1(G387), .A2(new_n1156), .A3(new_n1072), .A4(G375), .ZN(G407));
  NAND3_X1  g0957(.A1(new_n612), .A2(new_n613), .A3(G213), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(G375), .A2(new_n1072), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT122), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(G407), .A2(G213), .A3(new_n1160), .ZN(G409));
  INV_X1    g0961(.A(new_n1158), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1074), .A2(new_n1075), .A3(new_n1128), .A4(new_n1101), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1072), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT123), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1128), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1092), .A2(new_n1133), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1128), .A2(new_n1165), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1162), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT60), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1132), .B1(new_n1172), .B2(new_n1021), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1130), .A2(new_n1091), .A3(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(new_n637), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1152), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(G384), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(G384), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT63), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1171), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(G390), .A2(new_n915), .A3(new_n940), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G390), .B1(new_n915), .B2(new_n940), .ZN(new_n1185));
  OAI21_X1  g0985(.A(G396), .B1(new_n943), .B2(new_n976), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT126), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1155), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1155), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1184), .A2(new_n1185), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G387), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1189), .B1(new_n1192), .B2(new_n1183), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1182), .A2(new_n1194), .A3(KEYINPUT61), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT124), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1179), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT124), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1163), .A2(new_n1170), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1158), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1180), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1158), .A3(new_n1200), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G2897), .B(new_n1162), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1162), .A2(G2897), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1203), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1195), .A2(new_n1202), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT61), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n1171), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1215));
  NAND2_X1  g1015(.A1(new_n1201), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1171), .A2(KEYINPUT62), .A3(new_n1198), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1194), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1211), .B1(new_n1218), .B2(new_n1219), .ZN(G405));
  NAND2_X1  g1020(.A1(G375), .A2(new_n1164), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1163), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(new_n1198), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(new_n1194), .ZN(G402));
endmodule


