

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  XNOR2_X1 U326 ( .A(n452), .B(n451), .ZN(n458) );
  XNOR2_X1 U327 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U328 ( .A(n371), .B(n370), .Z(n577) );
  XOR2_X1 U329 ( .A(n358), .B(n357), .Z(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT119), .B(KEYINPUT45), .ZN(n337) );
  XNOR2_X1 U331 ( .A(KEYINPUT118), .B(KEYINPUT47), .ZN(n377) );
  XNOR2_X1 U332 ( .A(n338), .B(n337), .ZN(n373) );
  INV_X1 U333 ( .A(KEYINPUT102), .ZN(n471) );
  XNOR2_X1 U334 ( .A(n378), .B(n377), .ZN(n379) );
  INV_X1 U335 ( .A(n396), .ZN(n321) );
  XNOR2_X1 U336 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U337 ( .A(n479), .B(KEYINPUT104), .ZN(n480) );
  XNOR2_X1 U338 ( .A(n324), .B(n323), .ZN(n328) );
  XNOR2_X1 U339 ( .A(n481), .B(n480), .ZN(n533) );
  XNOR2_X1 U340 ( .A(n425), .B(KEYINPUT64), .ZN(n489) );
  INV_X1 U341 ( .A(KEYINPUT60), .ZN(n463) );
  XNOR2_X1 U342 ( .A(n492), .B(KEYINPUT123), .ZN(n582) );
  XOR2_X1 U343 ( .A(n336), .B(n335), .Z(n581) );
  XOR2_X1 U344 ( .A(n460), .B(n459), .Z(n524) );
  XNOR2_X1 U345 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U346 ( .A(n485), .B(G43GAT), .ZN(n486) );
  XNOR2_X1 U347 ( .A(n466), .B(n465), .ZN(G1352GAT) );
  XNOR2_X1 U348 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  INV_X1 U349 ( .A(KEYINPUT48), .ZN(n382) );
  XOR2_X1 U350 ( .A(G155GAT), .B(G211GAT), .Z(n296) );
  XNOR2_X1 U351 ( .A(G183GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(n297), .B(G78GAT), .Z(n299) );
  XOR2_X1 U354 ( .A(G1GAT), .B(KEYINPUT73), .Z(n363) );
  XNOR2_X1 U355 ( .A(G22GAT), .B(n363), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(G8GAT), .B(KEYINPUT82), .Z(n391) );
  XOR2_X1 U358 ( .A(n300), .B(n391), .Z(n303) );
  XOR2_X1 U359 ( .A(G15GAT), .B(G127GAT), .Z(n454) );
  XNOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT75), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n301), .B(KEYINPUT13), .ZN(n341) );
  XNOR2_X1 U362 ( .A(n454), .B(n341), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U364 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n305) );
  NAND2_X1 U365 ( .A1(G231GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U367 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U368 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n309) );
  XNOR2_X1 U369 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n310), .B(G64GAT), .ZN(n311) );
  XOR2_X1 U372 ( .A(n312), .B(n311), .Z(n572) );
  INV_X1 U373 ( .A(n572), .ZN(n588) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(KEYINPUT77), .ZN(n343) );
  INV_X1 U376 ( .A(n343), .ZN(n315) );
  INV_X1 U377 ( .A(G92GAT), .ZN(n314) );
  NAND2_X1 U378 ( .A1(n315), .A2(n314), .ZN(n317) );
  NAND2_X1 U379 ( .A1(n343), .A2(G92GAT), .ZN(n316) );
  NAND2_X1 U380 ( .A1(n317), .A2(n316), .ZN(n319) );
  AND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XOR2_X1 U384 ( .A(G134GAT), .B(KEYINPUT80), .Z(n416) );
  XNOR2_X1 U385 ( .A(n437), .B(n416), .ZN(n322) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n320), .B(KEYINPUT81), .ZN(n396) );
  XOR2_X1 U388 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n326) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U391 ( .A(n328), .B(n327), .Z(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT7), .B(KEYINPUT72), .Z(n330) );
  XNOR2_X1 U393 ( .A(G43GAT), .B(G29GAT), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U395 ( .A(KEYINPUT8), .B(n331), .Z(n370) );
  XOR2_X1 U396 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n333) );
  XNOR2_X1 U397 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n370), .B(n334), .ZN(n335) );
  XNOR2_X1 U400 ( .A(KEYINPUT36), .B(n581), .ZN(n590) );
  NAND2_X1 U401 ( .A1(n588), .A2(n590), .ZN(n338) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n392) );
  XOR2_X1 U405 ( .A(n392), .B(n341), .Z(n345) );
  XNOR2_X1 U406 ( .A(G106GAT), .B(G78GAT), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n342), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U408 ( .A(n430), .B(n343), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n352) );
  XOR2_X1 U410 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XOR2_X1 U411 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n347) );
  XNOR2_X1 U412 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U414 ( .A(n445), .B(n348), .Z(n350) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n482) );
  XOR2_X1 U418 ( .A(KEYINPUT69), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U419 ( .A(G113GAT), .B(G197GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U421 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n356) );
  XNOR2_X1 U422 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U424 ( .A(KEYINPUT30), .B(KEYINPUT74), .Z(n360) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT29), .B(n361), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n294), .B(n362), .ZN(n367) );
  XOR2_X1 U429 ( .A(G36GAT), .B(G50GAT), .Z(n365) );
  XOR2_X1 U430 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XNOR2_X1 U431 ( .A(n438), .B(n363), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U433 ( .A(n367), .B(n366), .Z(n369) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(G15GAT), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n371) );
  INV_X1 U436 ( .A(n577), .ZN(n565) );
  AND2_X1 U437 ( .A1(n482), .A2(n565), .ZN(n372) );
  AND2_X1 U438 ( .A1(n373), .A2(n372), .ZN(n380) );
  XOR2_X1 U439 ( .A(n482), .B(KEYINPUT41), .Z(n568) );
  NOR2_X1 U440 ( .A1(n565), .A2(n568), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n374), .B(KEYINPUT46), .ZN(n375) );
  NOR2_X1 U442 ( .A1(n588), .A2(n375), .ZN(n376) );
  INV_X1 U443 ( .A(n581), .ZN(n575) );
  NAND2_X1 U444 ( .A1(n376), .A2(n575), .ZN(n378) );
  NOR2_X1 U445 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n547) );
  XOR2_X1 U447 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT89), .B(KEYINPUT18), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U450 ( .A(n385), .B(KEYINPUT90), .Z(n387) );
  XNOR2_X1 U451 ( .A(G169GAT), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n452) );
  XOR2_X1 U453 ( .A(KEYINPUT94), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U454 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U456 ( .A(G197GAT), .B(n390), .Z(n442) );
  XNOR2_X1 U457 ( .A(n452), .B(n442), .ZN(n400) );
  XOR2_X1 U458 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U461 ( .A(n395), .B(KEYINPUT100), .Z(n398) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT101), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U464 ( .A(n400), .B(n399), .Z(n537) );
  XNOR2_X1 U465 ( .A(n537), .B(KEYINPUT122), .ZN(n401) );
  AND2_X1 U466 ( .A1(n547), .A2(n401), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT54), .ZN(n424) );
  XOR2_X1 U468 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n404) );
  XNOR2_X1 U469 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n423) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G120GAT), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U474 ( .A(G57GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(G127GAT), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U477 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n412) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U481 ( .A(G1GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U483 ( .A(n417), .B(n416), .Z(n421) );
  XOR2_X1 U484 ( .A(G113GAT), .B(KEYINPUT0), .Z(n453) );
  XOR2_X1 U485 ( .A(G155GAT), .B(KEYINPUT3), .Z(n419) );
  XNOR2_X1 U486 ( .A(KEYINPUT95), .B(KEYINPUT2), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n453), .B(n429), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U490 ( .A(n423), .B(n422), .Z(n535) );
  INV_X1 U491 ( .A(n535), .ZN(n518) );
  NAND2_X1 U492 ( .A1(n424), .A2(n518), .ZN(n425) );
  XOR2_X1 U493 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n427) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U496 ( .A(n428), .B(KEYINPUT93), .Z(n432) );
  XNOR2_X1 U497 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U499 ( .A(G204GAT), .B(KEYINPUT24), .Z(n434) );
  XNOR2_X1 U500 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U502 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n488) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT92), .Z(n444) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U509 ( .A(n446), .B(n445), .Z(n450) );
  XOR2_X1 U510 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n448) );
  XNOR2_X1 U511 ( .A(KEYINPUT88), .B(KEYINPUT91), .ZN(n447) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U513 ( .A(G190GAT), .B(G99GAT), .Z(n456) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U516 ( .A(n458), .B(n457), .Z(n460) );
  XNOR2_X1 U517 ( .A(G43GAT), .B(G134GAT), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n488), .A2(n524), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT26), .ZN(n563) );
  NOR2_X1 U520 ( .A1(n489), .A2(n563), .ZN(n591) );
  NAND2_X1 U521 ( .A1(n591), .A2(n577), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT59), .ZN(n466) );
  XNOR2_X1 U523 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n464) );
  XOR2_X1 U524 ( .A(n537), .B(KEYINPUT27), .Z(n474) );
  NOR2_X1 U525 ( .A1(n563), .A2(n474), .ZN(n470) );
  INV_X1 U526 ( .A(n537), .ZN(n522) );
  NOR2_X1 U527 ( .A1(n522), .A2(n524), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n488), .A2(n467), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NOR2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n518), .ZN(n477) );
  OR2_X1 U533 ( .A1(n518), .A2(n474), .ZN(n562) );
  XNOR2_X1 U534 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n475) );
  XOR2_X1 U535 ( .A(n475), .B(n488), .Z(n528) );
  INV_X1 U536 ( .A(n528), .ZN(n542) );
  NOR2_X1 U537 ( .A1(n562), .A2(n542), .ZN(n548) );
  NAND2_X1 U538 ( .A1(n548), .A2(n524), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n477), .A2(n476), .ZN(n499) );
  NAND2_X1 U540 ( .A1(n590), .A2(n499), .ZN(n478) );
  NOR2_X1 U541 ( .A1(n588), .A2(n478), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT105), .B(KEYINPUT37), .ZN(n479) );
  INV_X1 U543 ( .A(n482), .ZN(n585) );
  NOR2_X1 U544 ( .A1(n585), .A2(n565), .ZN(n501) );
  NAND2_X1 U545 ( .A1(n533), .A2(n501), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n483), .B(KEYINPUT38), .ZN(n484) );
  XNOR2_X1 U547 ( .A(KEYINPUT106), .B(n484), .ZN(n513) );
  NOR2_X1 U548 ( .A1(n513), .A2(n524), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n485) );
  NOR2_X1 U550 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT55), .B(n490), .Z(n491) );
  INV_X1 U552 ( .A(n524), .ZN(n549) );
  NAND2_X1 U553 ( .A1(n491), .A2(n549), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT108), .B(n568), .Z(n553) );
  NAND2_X1 U555 ( .A1(n582), .A2(n553), .ZN(n496) );
  XOR2_X1 U556 ( .A(G176GAT), .B(KEYINPUT56), .Z(n494) );
  XNOR2_X1 U557 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1349GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT86), .B(KEYINPUT16), .Z(n498) );
  NAND2_X1 U561 ( .A1(n588), .A2(n575), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n500) );
  AND2_X1 U563 ( .A1(n500), .A2(n499), .ZN(n516) );
  NAND2_X1 U564 ( .A1(n501), .A2(n516), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n518), .A2(n507), .ZN(n502) );
  XOR2_X1 U566 ( .A(G1GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT34), .B(n503), .ZN(G1324GAT) );
  NOR2_X1 U568 ( .A1(n522), .A2(n507), .ZN(n504) );
  XOR2_X1 U569 ( .A(G8GAT), .B(n504), .Z(G1325GAT) );
  NOR2_X1 U570 ( .A1(n524), .A2(n507), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  NOR2_X1 U573 ( .A1(n528), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  NOR2_X1 U576 ( .A1(n518), .A2(n513), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U579 ( .A1(n522), .A2(n513), .ZN(n512) );
  XOR2_X1 U580 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U581 ( .A1(n528), .A2(n513), .ZN(n514) );
  XOR2_X1 U582 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  NAND2_X1 U583 ( .A1(n553), .A2(n565), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(KEYINPUT109), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n532), .A2(n516), .ZN(n517) );
  XNOR2_X1 U586 ( .A(KEYINPUT110), .B(n517), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n527), .A2(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U590 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U591 ( .A1(n522), .A2(n527), .ZN(n523) );
  XOR2_X1 U592 ( .A(G64GAT), .B(n523), .Z(G1333GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n524), .ZN(n525) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(n525), .Z(n526) );
  XNOR2_X1 U595 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  XNOR2_X1 U596 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n530) );
  NOR2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(G78GAT), .B(n531), .Z(G1335GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(n534), .Z(n543) );
  NAND2_X1 U602 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U604 ( .A(G92GAT), .B(KEYINPUT115), .Z(n539) );
  NAND2_X1 U605 ( .A1(n543), .A2(n537), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1337GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n549), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(KEYINPUT116), .ZN(n541) );
  XNOR2_X1 U609 ( .A(G99GAT), .B(n541), .ZN(G1338GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT44), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  INV_X1 U614 ( .A(n547), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n559), .A2(n577), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U619 ( .A(G120GAT), .B(KEYINPUT49), .Z(n555) );
  NAND2_X1 U620 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1341GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n557) );
  NAND2_X1 U623 ( .A1(n559), .A2(n588), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G127GAT), .B(n558), .Z(G1342GAT) );
  XOR2_X1 U626 ( .A(G134GAT), .B(KEYINPUT51), .Z(n561) );
  NAND2_X1 U627 ( .A1(n559), .A2(n581), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1343GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n547), .A2(n564), .ZN(n574) );
  NOR2_X1 U631 ( .A1(n565), .A2(n574), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1344GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n574), .ZN(n570) );
  XNOR2_X1 U635 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G148GAT), .B(n571), .ZN(G1345GAT) );
  NOR2_X1 U638 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U639 ( .A(G155GAT), .B(n573), .Z(G1346GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G162GAT), .B(n576), .Z(G1347GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n582), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G169GAT), .B(n578), .ZN(G1348GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U645 ( .A1(n582), .A2(n588), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1350GAT) );
  XNOR2_X1 U647 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1351GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n591), .A2(n588), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n593) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

