

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n520), .ZN(n725) );
  BUF_X2 U556 ( .A(n749), .Z(n520) );
  XNOR2_X1 U557 ( .A(n698), .B(KEYINPUT64), .ZN(n749) );
  INV_X1 U558 ( .A(n548), .ZN(n563) );
  XNOR2_X1 U559 ( .A(n758), .B(n757), .ZN(n774) );
  XOR2_X1 U560 ( .A(KEYINPUT72), .B(n593), .Z(n992) );
  NOR2_X2 U561 ( .A1(G2104), .A2(n552), .ZN(n901) );
  BUF_X2 U562 ( .A(n804), .Z(n521) );
  NOR2_X1 U563 ( .A1(G1961), .A2(n725), .ZN(n724) );
  NOR2_X1 U564 ( .A1(G171), .A2(n736), .ZN(n737) );
  INV_X1 U565 ( .A(KEYINPUT65), .ZN(n764) );
  AND2_X1 U566 ( .A1(n827), .A2(n821), .ZN(n815) );
  NOR2_X1 U567 ( .A1(n733), .A2(G168), .ZN(n735) );
  NAND2_X1 U568 ( .A1(n742), .A2(n741), .ZN(n748) );
  XNOR2_X1 U569 ( .A(n740), .B(KEYINPUT31), .ZN(n741) );
  INV_X1 U570 ( .A(KEYINPUT33), .ZN(n767) );
  INV_X1 U571 ( .A(n977), .ZN(n770) );
  INV_X1 U572 ( .A(KEYINPUT106), .ZN(n817) );
  OR2_X1 U573 ( .A1(n784), .A2(n783), .ZN(n522) );
  NOR2_X1 U574 ( .A1(n771), .A2(n770), .ZN(n523) );
  NOR2_X1 U575 ( .A1(n745), .A2(n744), .ZN(n524) );
  AND2_X1 U576 ( .A1(n780), .A2(n779), .ZN(n525) );
  NOR2_X1 U577 ( .A1(n520), .A2(n956), .ZN(n699) );
  NOR2_X1 U578 ( .A1(n702), .A2(n992), .ZN(n709) );
  NOR2_X1 U579 ( .A1(n715), .A2(n714), .ZN(n718) );
  INV_X1 U580 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U581 ( .A(n723), .B(n722), .ZN(n729) );
  INV_X1 U582 ( .A(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U583 ( .A1(n748), .A2(n524), .ZN(n773) );
  NOR2_X1 U584 ( .A1(n695), .A2(G1384), .ZN(n696) );
  INV_X1 U585 ( .A(KEYINPUT17), .ZN(n546) );
  XNOR2_X1 U586 ( .A(n697), .B(KEYINPUT95), .ZN(n786) );
  INV_X1 U587 ( .A(n786), .ZN(n787) );
  XNOR2_X1 U588 ( .A(n818), .B(n817), .ZN(n820) );
  NOR2_X2 U589 ( .A1(G651), .A2(G543), .ZN(n657) );
  NOR2_X1 U590 ( .A1(G651), .A2(n647), .ZN(n661) );
  XNOR2_X1 U591 ( .A(n576), .B(KEYINPUT91), .ZN(n577) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n647) );
  NAND2_X1 U593 ( .A1(G52), .A2(n661), .ZN(n528) );
  INV_X1 U594 ( .A(G651), .ZN(n529) );
  NOR2_X1 U595 ( .A1(G543), .A2(n529), .ZN(n526) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n526), .Z(n662) );
  NAND2_X1 U597 ( .A1(G64), .A2(n662), .ZN(n527) );
  NAND2_X1 U598 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U599 ( .A1(G90), .A2(n657), .ZN(n531) );
  NOR2_X1 U600 ( .A1(n647), .A2(n529), .ZN(n658) );
  NAND2_X1 U601 ( .A1(G77), .A2(n658), .ZN(n530) );
  NAND2_X1 U602 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n532), .Z(n533) );
  NOR2_X1 U604 ( .A1(n534), .A2(n533), .ZN(G171) );
  NAND2_X1 U605 ( .A1(G51), .A2(n661), .ZN(n536) );
  NAND2_X1 U606 ( .A1(G63), .A2(n662), .ZN(n535) );
  NAND2_X1 U607 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U608 ( .A(KEYINPUT6), .B(n537), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n657), .A2(G89), .ZN(n538) );
  XNOR2_X1 U610 ( .A(n538), .B(KEYINPUT4), .ZN(n540) );
  NAND2_X1 U611 ( .A1(G76), .A2(n658), .ZN(n539) );
  NAND2_X1 U612 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U613 ( .A(n541), .B(KEYINPUT5), .Z(n542) );
  NOR2_X1 U614 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(n544), .Z(n545) );
  XNOR2_X1 U616 ( .A(KEYINPUT76), .B(n545), .ZN(G168) );
  NOR2_X1 U617 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n547), .B(n546), .ZN(n568) );
  INV_X1 U619 ( .A(n568), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n563), .A2(G137), .ZN(n551) );
  INV_X1 U621 ( .A(G2104), .ZN(n553) );
  NOR2_X1 U622 ( .A1(G2105), .A2(n553), .ZN(n804) );
  NAND2_X1 U623 ( .A1(G101), .A2(n804), .ZN(n549) );
  XOR2_X1 U624 ( .A(KEYINPUT23), .B(n549), .Z(n550) );
  NAND2_X1 U625 ( .A1(n551), .A2(n550), .ZN(n557) );
  INV_X1 U626 ( .A(G2105), .ZN(n552) );
  NOR2_X1 U627 ( .A1(n553), .A2(n552), .ZN(n572) );
  BUF_X1 U628 ( .A(n572), .Z(n900) );
  NAND2_X1 U629 ( .A1(G113), .A2(n900), .ZN(n555) );
  NAND2_X1 U630 ( .A1(G125), .A2(n901), .ZN(n554) );
  NAND2_X1 U631 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U632 ( .A1(n557), .A2(n556), .ZN(G160) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U634 ( .A1(G111), .A2(n900), .ZN(n559) );
  NAND2_X1 U635 ( .A1(G99), .A2(n521), .ZN(n558) );
  NAND2_X1 U636 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U637 ( .A1(n901), .A2(G123), .ZN(n560) );
  XOR2_X1 U638 ( .A(KEYINPUT18), .B(n560), .Z(n561) );
  NOR2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n563), .A2(G135), .ZN(n564) );
  NAND2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n939) );
  XNOR2_X1 U642 ( .A(G2096), .B(n939), .ZN(n566) );
  OR2_X1 U643 ( .A1(G2100), .A2(n566), .ZN(G156) );
  NAND2_X1 U644 ( .A1(G102), .A2(n521), .ZN(n567) );
  XNOR2_X1 U645 ( .A(n567), .B(KEYINPUT92), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n568), .A2(G138), .ZN(n569) );
  XOR2_X1 U647 ( .A(n569), .B(KEYINPUT93), .Z(n570) );
  NAND2_X1 U648 ( .A1(n571), .A2(n570), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n572), .A2(G114), .ZN(n573) );
  XNOR2_X1 U650 ( .A(n573), .B(KEYINPUT90), .ZN(n575) );
  NAND2_X1 U651 ( .A1(G126), .A2(n901), .ZN(n574) );
  AND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n695) );
  BUF_X1 U654 ( .A(n695), .Z(G164) );
  INV_X1 U655 ( .A(G82), .ZN(G220) );
  INV_X1 U656 ( .A(G120), .ZN(G236) );
  INV_X1 U657 ( .A(G69), .ZN(G235) );
  INV_X1 U658 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U659 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n579) );
  XNOR2_X1 U660 ( .A(n579), .B(G168), .ZN(G286) );
  XOR2_X1 U661 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n581) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U663 ( .A(n581), .B(n580), .ZN(G223) );
  XOR2_X1 U664 ( .A(G223), .B(KEYINPUT70), .Z(n839) );
  NAND2_X1 U665 ( .A1(n839), .A2(G567), .ZN(n582) );
  XOR2_X1 U666 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  XOR2_X1 U667 ( .A(G860), .B(KEYINPUT73), .Z(n615) );
  NAND2_X1 U668 ( .A1(G81), .A2(n657), .ZN(n583) );
  XOR2_X1 U669 ( .A(KEYINPUT71), .B(n583), .Z(n584) );
  XNOR2_X1 U670 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U671 ( .A1(G68), .A2(n658), .ZN(n585) );
  NAND2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U673 ( .A(n587), .B(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U674 ( .A1(G43), .A2(n661), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U676 ( .A1(n662), .A2(G56), .ZN(n590) );
  XOR2_X1 U677 ( .A(KEYINPUT14), .B(n590), .Z(n591) );
  NOR2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U679 ( .A(n992), .ZN(n594) );
  NAND2_X1 U680 ( .A1(n615), .A2(n594), .ZN(G153) );
  INV_X1 U681 ( .A(G171), .ZN(G301) );
  NAND2_X1 U682 ( .A1(G66), .A2(n662), .ZN(n601) );
  NAND2_X1 U683 ( .A1(G79), .A2(n658), .ZN(n596) );
  NAND2_X1 U684 ( .A1(G54), .A2(n661), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U686 ( .A1(n657), .A2(G92), .ZN(n597) );
  XOR2_X1 U687 ( .A(KEYINPUT74), .B(n597), .Z(n598) );
  NOR2_X1 U688 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U690 ( .A(n602), .B(KEYINPUT15), .ZN(n916) );
  NOR2_X1 U691 ( .A1(n916), .A2(G868), .ZN(n603) );
  XNOR2_X1 U692 ( .A(n603), .B(KEYINPUT75), .ZN(n605) );
  NAND2_X1 U693 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U695 ( .A1(G53), .A2(n661), .ZN(n607) );
  NAND2_X1 U696 ( .A1(G65), .A2(n662), .ZN(n606) );
  NAND2_X1 U697 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U698 ( .A1(G91), .A2(n657), .ZN(n609) );
  NAND2_X1 U699 ( .A1(G78), .A2(n658), .ZN(n608) );
  NAND2_X1 U700 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U701 ( .A1(n611), .A2(n610), .ZN(n980) );
  INV_X1 U702 ( .A(n980), .ZN(G299) );
  NAND2_X1 U703 ( .A1(G868), .A2(G286), .ZN(n613) );
  INV_X1 U704 ( .A(G868), .ZN(n677) );
  NAND2_X1 U705 ( .A1(G299), .A2(n677), .ZN(n612) );
  NAND2_X1 U706 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U707 ( .A(n916), .ZN(n982) );
  INV_X1 U708 ( .A(G559), .ZN(n614) );
  NOR2_X1 U709 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U710 ( .A1(n982), .A2(n616), .ZN(n617) );
  XOR2_X1 U711 ( .A(n617), .B(KEYINPUT16), .Z(n618) );
  XNOR2_X1 U712 ( .A(KEYINPUT78), .B(n618), .ZN(G148) );
  NOR2_X1 U713 ( .A1(G559), .A2(n677), .ZN(n619) );
  NAND2_X1 U714 ( .A1(n916), .A2(n619), .ZN(n620) );
  XNOR2_X1 U715 ( .A(n620), .B(KEYINPUT79), .ZN(n622) );
  NOR2_X1 U716 ( .A1(n992), .A2(G868), .ZN(n621) );
  NOR2_X1 U717 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U718 ( .A1(G559), .A2(n916), .ZN(n623) );
  XNOR2_X1 U719 ( .A(n623), .B(KEYINPUT80), .ZN(n675) );
  XOR2_X1 U720 ( .A(n992), .B(n675), .Z(n624) );
  XNOR2_X1 U721 ( .A(KEYINPUT81), .B(n624), .ZN(n625) );
  NOR2_X1 U722 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U723 ( .A(n626), .B(KEYINPUT82), .Z(n634) );
  NAND2_X1 U724 ( .A1(G93), .A2(n657), .ZN(n628) );
  NAND2_X1 U725 ( .A1(G80), .A2(n658), .ZN(n627) );
  NAND2_X1 U726 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U727 ( .A1(G55), .A2(n661), .ZN(n629) );
  XNOR2_X1 U728 ( .A(KEYINPUT83), .B(n629), .ZN(n630) );
  NOR2_X1 U729 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U730 ( .A1(n662), .A2(G67), .ZN(n632) );
  NAND2_X1 U731 ( .A1(n633), .A2(n632), .ZN(n678) );
  XNOR2_X1 U732 ( .A(n634), .B(n678), .ZN(G145) );
  NAND2_X1 U733 ( .A1(G73), .A2(n658), .ZN(n635) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(n635), .Z(n640) );
  NAND2_X1 U735 ( .A1(G86), .A2(n657), .ZN(n637) );
  NAND2_X1 U736 ( .A1(G61), .A2(n662), .ZN(n636) );
  NAND2_X1 U737 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U738 ( .A(KEYINPUT85), .B(n638), .Z(n639) );
  NOR2_X1 U739 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U740 ( .A1(n661), .A2(G48), .ZN(n641) );
  NAND2_X1 U741 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U742 ( .A1(G49), .A2(n661), .ZN(n644) );
  NAND2_X1 U743 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U744 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U745 ( .A(KEYINPUT84), .B(n645), .ZN(n646) );
  NOR2_X1 U746 ( .A1(n662), .A2(n646), .ZN(n649) );
  NAND2_X1 U747 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U748 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U749 ( .A1(G85), .A2(n657), .ZN(n651) );
  NAND2_X1 U750 ( .A1(G72), .A2(n658), .ZN(n650) );
  NAND2_X1 U751 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U752 ( .A(KEYINPUT67), .B(n652), .ZN(n656) );
  NAND2_X1 U753 ( .A1(G47), .A2(n661), .ZN(n654) );
  NAND2_X1 U754 ( .A1(G60), .A2(n662), .ZN(n653) );
  AND2_X1 U755 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U756 ( .A1(n656), .A2(n655), .ZN(G290) );
  NAND2_X1 U757 ( .A1(G88), .A2(n657), .ZN(n660) );
  NAND2_X1 U758 ( .A1(G75), .A2(n658), .ZN(n659) );
  NAND2_X1 U759 ( .A1(n660), .A2(n659), .ZN(n666) );
  NAND2_X1 U760 ( .A1(G50), .A2(n661), .ZN(n664) );
  NAND2_X1 U761 ( .A1(G62), .A2(n662), .ZN(n663) );
  NAND2_X1 U762 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U763 ( .A1(n666), .A2(n665), .ZN(G166) );
  XNOR2_X1 U764 ( .A(G305), .B(G288), .ZN(n672) );
  XNOR2_X1 U765 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n668) );
  XNOR2_X1 U766 ( .A(G290), .B(G166), .ZN(n667) );
  XNOR2_X1 U767 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U768 ( .A(n980), .B(n669), .ZN(n670) );
  XNOR2_X1 U769 ( .A(n670), .B(n678), .ZN(n671) );
  XNOR2_X1 U770 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U771 ( .A(n992), .B(n673), .ZN(n915) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(n915), .ZN(n674) );
  XNOR2_X1 U773 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U774 ( .A1(n677), .A2(n676), .ZN(n680) );
  NOR2_X1 U775 ( .A1(G868), .A2(n678), .ZN(n679) );
  NOR2_X1 U776 ( .A1(n680), .A2(n679), .ZN(G295) );
  XOR2_X1 U777 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n682) );
  NAND2_X1 U778 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XNOR2_X1 U779 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U780 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U781 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U782 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U783 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U784 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U785 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U786 ( .A(n686), .B(KEYINPUT89), .ZN(n687) );
  NOR2_X1 U787 ( .A1(G238), .A2(n687), .ZN(n688) );
  NAND2_X1 U788 ( .A1(G57), .A2(n688), .ZN(n844) );
  NAND2_X1 U789 ( .A1(n844), .A2(G567), .ZN(n693) );
  NOR2_X1 U790 ( .A1(G219), .A2(G220), .ZN(n689) );
  XOR2_X1 U791 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U792 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U793 ( .A1(G96), .A2(n691), .ZN(n845) );
  NAND2_X1 U794 ( .A1(n845), .A2(G2106), .ZN(n692) );
  NAND2_X1 U795 ( .A1(n693), .A2(n692), .ZN(n926) );
  NAND2_X1 U796 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U797 ( .A1(n926), .A2(n694), .ZN(n843) );
  NAND2_X1 U798 ( .A1(n843), .A2(G36), .ZN(G176) );
  XOR2_X1 U799 ( .A(KEYINPUT94), .B(G166), .Z(G303) );
  XNOR2_X1 U800 ( .A(n696), .B(KEYINPUT66), .ZN(n785) );
  NAND2_X1 U801 ( .A1(G40), .A2(G160), .ZN(n697) );
  NAND2_X1 U802 ( .A1(n785), .A2(n786), .ZN(n698) );
  INV_X1 U803 ( .A(G1996), .ZN(n956) );
  XOR2_X1 U804 ( .A(n699), .B(KEYINPUT26), .Z(n701) );
  NAND2_X1 U805 ( .A1(n520), .A2(G1341), .ZN(n700) );
  NAND2_X1 U806 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U807 ( .A1(n709), .A2(n916), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n520), .A2(G1348), .ZN(n703) );
  XNOR2_X1 U809 ( .A(n703), .B(KEYINPUT102), .ZN(n705) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n725), .ZN(n704) );
  NAND2_X1 U811 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U812 ( .A(KEYINPUT103), .B(n706), .Z(n707) );
  NAND2_X1 U813 ( .A1(n708), .A2(n707), .ZN(n711) );
  OR2_X1 U814 ( .A1(n916), .A2(n709), .ZN(n710) );
  NAND2_X1 U815 ( .A1(n711), .A2(n710), .ZN(n717) );
  NAND2_X1 U816 ( .A1(G2072), .A2(n725), .ZN(n712) );
  XNOR2_X1 U817 ( .A(KEYINPUT27), .B(n712), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n520), .A2(G1956), .ZN(n713) );
  XNOR2_X1 U819 ( .A(KEYINPUT101), .B(n713), .ZN(n714) );
  NAND2_X1 U820 ( .A1(n718), .A2(n980), .ZN(n716) );
  NAND2_X1 U821 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U822 ( .A1(n718), .A2(n980), .ZN(n719) );
  XOR2_X1 U823 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U824 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U825 ( .A(KEYINPUT100), .B(n724), .Z(n727) );
  XNOR2_X1 U826 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U827 ( .A1(n725), .A2(n955), .ZN(n726) );
  NAND2_X1 U828 ( .A1(n727), .A2(n726), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G171), .ZN(n728) );
  NAND2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n520), .A2(G8), .ZN(n784) );
  NOR2_X1 U832 ( .A1(G1966), .A2(n784), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n520), .A2(G2084), .ZN(n743) );
  INV_X1 U834 ( .A(n743), .ZN(n730) );
  NAND2_X1 U835 ( .A1(n730), .A2(G8), .ZN(n731) );
  OR2_X1 U836 ( .A1(n744), .A2(n731), .ZN(n732) );
  XNOR2_X1 U837 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  INV_X1 U838 ( .A(KEYINPUT104), .ZN(n734) );
  XNOR2_X1 U839 ( .A(n735), .B(n734), .ZN(n739) );
  XNOR2_X1 U840 ( .A(KEYINPUT105), .B(n737), .ZN(n738) );
  NAND2_X1 U841 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U842 ( .A1(G8), .A2(n743), .ZN(n745) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U844 ( .A(n996), .ZN(n746) );
  OR2_X1 U845 ( .A1(n784), .A2(n746), .ZN(n761) );
  INV_X1 U846 ( .A(n761), .ZN(n747) );
  AND2_X1 U847 ( .A1(n773), .A2(n747), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n748), .A2(G286), .ZN(n756) );
  INV_X1 U849 ( .A(G8), .ZN(n754) );
  NOR2_X1 U850 ( .A1(G1971), .A2(n784), .ZN(n751) );
  NOR2_X1 U851 ( .A1(n520), .A2(G2090), .ZN(n750) );
  NOR2_X1 U852 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U853 ( .A1(n752), .A2(G303), .ZN(n753) );
  OR2_X1 U854 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U855 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U856 ( .A1(n759), .A2(n774), .ZN(n763) );
  NOR2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n995) );
  NOR2_X1 U858 ( .A1(G303), .A2(G1971), .ZN(n1002) );
  NOR2_X1 U859 ( .A1(n995), .A2(n1002), .ZN(n760) );
  OR2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U861 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U862 ( .A(n765), .B(n764), .ZN(n766) );
  INV_X1 U863 ( .A(n766), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n995), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U866 ( .A1(n769), .A2(n784), .ZN(n771) );
  XOR2_X1 U867 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U868 ( .A1(n772), .A2(n523), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n777) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U871 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n778), .A2(n784), .ZN(n779) );
  NOR2_X1 U874 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XNOR2_X1 U875 ( .A(n781), .B(KEYINPUT24), .ZN(n782) );
  XNOR2_X1 U876 ( .A(n782), .B(KEYINPUT99), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n525), .A2(n522), .ZN(n816) );
  NOR2_X1 U878 ( .A1(n785), .A2(n787), .ZN(n833) );
  NAND2_X1 U879 ( .A1(G104), .A2(n521), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G140), .A2(n563), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U882 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G116), .A2(n900), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G128), .A2(n901), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U888 ( .A(KEYINPUT36), .B(n796), .Z(n911) );
  XOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .Z(n829) );
  AND2_X1 U890 ( .A1(n911), .A2(n829), .ZN(n946) );
  NAND2_X1 U891 ( .A1(n833), .A2(n946), .ZN(n827) );
  NAND2_X1 U892 ( .A1(G107), .A2(n900), .ZN(n798) );
  NAND2_X1 U893 ( .A1(G95), .A2(n521), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n563), .A2(G131), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT96), .B(n799), .Z(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n901), .A2(G119), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n896) );
  AND2_X1 U900 ( .A1(n896), .A2(G1991), .ZN(n938) );
  NAND2_X1 U901 ( .A1(G105), .A2(n521), .ZN(n805) );
  XNOR2_X1 U902 ( .A(n805), .B(KEYINPUT38), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G117), .A2(n900), .ZN(n807) );
  NAND2_X1 U904 ( .A1(G129), .A2(n901), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U906 ( .A1(G141), .A2(n563), .ZN(n808) );
  XNOR2_X1 U907 ( .A(KEYINPUT97), .B(n808), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U910 ( .A(KEYINPUT98), .B(n813), .Z(n897) );
  NOR2_X1 U911 ( .A1(n956), .A2(n897), .ZN(n942) );
  OR2_X1 U912 ( .A1(n938), .A2(n942), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n833), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U915 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U916 ( .A1(n984), .A2(n833), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n836) );
  AND2_X1 U918 ( .A1(n956), .A2(n897), .ZN(n933) );
  INV_X1 U919 ( .A(n821), .ZN(n824) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n896), .ZN(n937) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n937), .A2(n822), .ZN(n823) );
  NOR2_X1 U923 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U924 ( .A1(n933), .A2(n825), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n826), .B(KEYINPUT39), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n829), .A2(n911), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(KEYINPUT107), .ZN(n947) );
  NAND2_X1 U929 ( .A1(n831), .A2(n947), .ZN(n832) );
  XNOR2_X1 U930 ( .A(KEYINPUT108), .B(n832), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(G329) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n839), .ZN(G217) );
  NAND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(n840), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n841), .A2(G661), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G188) );
  NOR2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G325) );
  XOR2_X1 U942 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U945 ( .A(G1348), .B(G2454), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n846), .B(G2430), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n847), .B(G1341), .ZN(n853) );
  XOR2_X1 U948 ( .A(G2443), .B(G2427), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2438), .B(G2446), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U951 ( .A(G2451), .B(G2435), .Z(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n854), .A2(G14), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(n855), .Z(G401) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2072), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2078), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n858), .B(G2096), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2090), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U962 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n862) );
  XNOR2_X1 U963 ( .A(G2678), .B(G2100), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(G227) );
  XNOR2_X1 U966 ( .A(G1956), .B(KEYINPUT41), .ZN(n874) );
  XOR2_X1 U967 ( .A(G1976), .B(G1981), .Z(n866) );
  XNOR2_X1 U968 ( .A(G1966), .B(G1971), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U970 ( .A(G1961), .B(G1986), .Z(n868) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U973 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U974 ( .A(G2474), .B(KEYINPUT114), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G124), .A2(n901), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n900), .A2(G112), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G100), .A2(n521), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G136), .A2(n563), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U984 ( .A1(n881), .A2(n880), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n883) );
  XNOR2_X1 U986 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U987 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n939), .B(n884), .ZN(n886) );
  XNOR2_X1 U989 ( .A(G160), .B(G162), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G115), .A2(n900), .ZN(n888) );
  NAND2_X1 U992 ( .A1(G127), .A2(n901), .ZN(n887) );
  NAND2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U994 ( .A(n889), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U995 ( .A1(G103), .A2(n521), .ZN(n890) );
  NAND2_X1 U996 ( .A1(n891), .A2(n890), .ZN(n894) );
  NAND2_X1 U997 ( .A1(n563), .A2(G139), .ZN(n892) );
  XOR2_X1 U998 ( .A(KEYINPUT116), .B(n892), .Z(n893) );
  NOR2_X1 U999 ( .A1(n894), .A2(n893), .ZN(n927) );
  XOR2_X1 U1000 ( .A(n895), .B(n927), .Z(n899) );
  XNOR2_X1 U1001 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(n899), .B(n898), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n900), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(G130), .A2(n901), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G106), .A2(n521), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(G142), .A2(n563), .ZN(n904) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1009 ( .A(KEYINPUT45), .B(n906), .Z(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1011 ( .A(n910), .B(n909), .Z(n913) );
  XNOR2_X1 U1012 ( .A(G164), .B(n911), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n914), .ZN(G395) );
  XOR2_X1 U1015 ( .A(KEYINPUT118), .B(n915), .Z(n918) );
  XNOR2_X1 U1016 ( .A(G171), .B(n916), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(n919), .B(G286), .Z(n920) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n920), .ZN(G397) );
  OR2_X1 U1020 ( .A1(n926), .A2(G401), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(n926), .ZN(G319) );
  INV_X1 U1028 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G164), .B(G2078), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(KEYINPUT50), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(n931), .B(KEYINPUT119), .ZN(n936) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n934), .Z(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n950) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n973), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n953), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n968) );
  XOR2_X1 U1051 ( .A(G25), .B(G1991), .Z(n954) );
  NAND2_X1 U1052 ( .A1(n954), .A2(G28), .ZN(n965) );
  XOR2_X1 U1053 ( .A(n955), .B(G27), .Z(n958) );
  XOR2_X1 U1054 ( .A(n956), .B(G32), .Z(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n959), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n966), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n969) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n969), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n973), .B(n972), .ZN(n975) );
  INV_X1 U1068 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n976), .ZN(n1036) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT57), .B(n979), .ZN(n991) );
  XNOR2_X1 U1075 ( .A(G1956), .B(n980), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT122), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1348), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1080 ( .A(G1961), .B(G301), .Z(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1005) );
  INV_X1 U1086 ( .A(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT123), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT124), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1034) );
  INV_X1 U1095 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1096 ( .A(KEYINPUT125), .B(G1961), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1008), .B(G5), .ZN(n1022) );
  XOR2_X1 U1098 ( .A(G1341), .B(G19), .Z(n1010) );
  XOR2_X1 U1099 ( .A(G1981), .B(G6), .Z(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1013), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT127), .B(G4), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1014) );
  XNOR2_X1 U1106 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT60), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G21), .B(G1966), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(G1971), .B(G22), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(G23), .B(G1976), .ZN(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XOR2_X1 U1115 ( .A(G1986), .B(G24), .Z(n1025) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(KEYINPUT58), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

