//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT64), .B(G50), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT65), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n254), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n257), .B1(G238), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n232), .A2(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G97), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT70), .B1(new_n268), .B2(new_n258), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n249), .A2(new_n250), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(new_n266), .C2(new_n267), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n260), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT71), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n260), .B(new_n275), .C1(new_n269), .C2(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(KEYINPUT13), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n260), .B(new_n278), .C1(new_n269), .C2(new_n272), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G190), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n216), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n207), .A2(KEYINPUT66), .A3(G33), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT66), .B1(new_n207), .B2(G33), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G77), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n283), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n283), .A2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n289), .B1(new_n206), .B2(G20), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n297), .A2(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n292), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n279), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(G200), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n280), .A2(new_n306), .A3(KEYINPUT72), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT72), .B1(new_n280), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT8), .B(G58), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n286), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n288), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n282), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT9), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n294), .A2(new_n207), .A3(G1), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n300), .A2(new_n317), .B1(new_n202), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n315), .B2(new_n319), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n256), .A2(new_n257), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n271), .B1(new_n329), .B2(new_n220), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G222), .A2(G1698), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n263), .A2(G223), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n261), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n330), .A2(new_n333), .B1(new_n259), .B2(G226), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT10), .B1(new_n323), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n322), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT69), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n320), .ZN(new_n342));
  INV_X1    g0142(.A(new_n335), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT10), .B1(new_n343), .B2(G190), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n344), .A3(new_n336), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n323), .A2(new_n341), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n335), .B1(new_n315), .B2(new_n319), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(G179), .B2(new_n335), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n256), .A2(new_n257), .B1(G244), .B2(new_n259), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n261), .A2(G232), .A3(new_n263), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n222), .B2(new_n261), .ZN(new_n354));
  INV_X1    g0154(.A(G238), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n329), .A2(new_n355), .A3(new_n263), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n258), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G200), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT67), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n286), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n311), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n283), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n206), .A2(G20), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n300), .A2(G77), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G77), .B2(new_n296), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n368), .A2(KEYINPUT68), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(KEYINPUT68), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n359), .B1(new_n337), .B2(new_n358), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n368), .ZN(new_n372));
  INV_X1    g0172(.A(G179), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n352), .A2(new_n357), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n358), .A2(new_n348), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n309), .A2(new_n351), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT75), .B1(new_n327), .B2(G33), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(new_n325), .A3(KEYINPUT3), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n381), .A3(new_n328), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n262), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G223), .B2(G1698), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n382), .A2(new_n384), .B1(new_n325), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n386), .A2(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n259), .A2(G232), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n254), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n255), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n387), .A2(new_n390), .A3(G179), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n258), .A2(new_n254), .A3(new_n232), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n256), .B2(new_n257), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n258), .ZN(new_n394));
  AOI21_X1  g0194(.A(G169), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT77), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n348), .B1(new_n387), .B2(new_n390), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n373), .A3(new_n394), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT77), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n382), .A2(new_n207), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n289), .B1(new_n402), .B2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n382), .A2(new_n404), .A3(new_n207), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G58), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n289), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n201), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT76), .B(G20), .C1(new_n408), .C2(new_n201), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(G159), .B2(new_n288), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n411), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  INV_X1    g0216(.A(G159), .ZN(new_n417));
  INV_X1    g0217(.A(new_n288), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n411), .B(new_n412), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n404), .B1(new_n261), .B2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n289), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n416), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n282), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n311), .A2(new_n365), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n299), .B1(new_n296), .B2(new_n311), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n401), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n396), .A2(new_n400), .B1(new_n424), .B2(new_n427), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n387), .A2(new_n390), .A3(new_n337), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n393), .B2(new_n394), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n424), .A2(new_n438), .A3(new_n427), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n424), .A2(new_n438), .A3(new_n441), .A4(new_n427), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n434), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n424), .A2(new_n438), .A3(new_n427), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(KEYINPUT17), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n433), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n279), .A2(G179), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n277), .A2(new_n447), .A3(KEYINPUT74), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT74), .B1(new_n277), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n305), .A2(G169), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n348), .B(new_n455), .C1(new_n304), .C2(new_n279), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n456), .B2(new_n453), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n303), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n378), .A2(new_n446), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n379), .A2(new_n381), .A3(G244), .A4(new_n328), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G1698), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n460), .A2(new_n221), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n261), .A2(new_n263), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n261), .A2(KEYINPUT80), .A3(new_n263), .A4(new_n463), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n462), .A2(new_n466), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n258), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G45), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n252), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n474), .B2(G41), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n478), .A4(new_n251), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n253), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(G41), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n478), .A2(new_n476), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n271), .ZN(new_n483));
  INV_X1    g0283(.A(G257), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n472), .A2(new_n373), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n492), .A2(new_n207), .B1(new_n220), .B2(new_n418), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n222), .B1(new_n420), .B2(new_n421), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n282), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n296), .B2(G97), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n318), .A2(KEYINPUT79), .A3(new_n489), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n283), .B(new_n296), .C1(G1), .C2(new_n325), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n489), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n485), .B1(new_n471), .B2(new_n258), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n487), .B(new_n502), .C1(G169), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n472), .A2(G190), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n491), .A2(new_n488), .ZN(new_n506));
  INV_X1    g0306(.A(new_n490), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n288), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n420), .A2(new_n421), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n500), .B1(new_n512), .B2(new_n282), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n505), .B(new_n513), .C1(new_n436), .C2(new_n503), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n355), .A2(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n379), .A2(new_n381), .A3(new_n328), .A4(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n461), .B2(new_n263), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n271), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  OR3_X1    g0322(.A1(new_n253), .A2(KEYINPUT82), .A3(G1), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n271), .A4(G250), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n251), .A2(new_n480), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT67), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n360), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n360), .A2(new_n529), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n296), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n499), .A2(new_n385), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n379), .A2(new_n381), .A3(new_n328), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(KEYINPUT84), .A3(new_n207), .A4(G68), .ZN(new_n535));
  NAND3_X1  g0335(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n207), .A2(new_n536), .B1(new_n537), .B2(new_n385), .ZN(new_n538));
  OAI21_X1  g0338(.A(G97), .B1(new_n284), .B2(new_n285), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n379), .A2(new_n381), .A3(new_n207), .A4(new_n328), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n289), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n535), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n532), .B(new_n533), .C1(new_n545), .C2(new_n282), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n327), .A2(KEYINPUT75), .A3(G33), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(KEYINPUT83), .A3(new_n379), .A4(new_n516), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n517), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n258), .B1(new_n553), .B2(new_n520), .ZN(new_n554));
  INV_X1    g0354(.A(new_n527), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(G190), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n528), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n348), .B1(new_n522), .B2(new_n527), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n545), .A2(new_n282), .ZN(new_n559));
  INV_X1    g0359(.A(new_n532), .ZN(new_n560));
  INV_X1    g0360(.A(new_n499), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n361), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n554), .A2(new_n373), .A3(new_n555), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n515), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n499), .A2(G116), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n296), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(G20), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n282), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n282), .A2(KEYINPUT86), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n468), .B(new_n207), .C1(G33), .C2(new_n489), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n282), .A2(KEYINPUT86), .A3(new_n572), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT86), .B1(new_n282), .B2(new_n572), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT20), .B(new_n578), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n571), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n223), .A2(new_n263), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n379), .A2(new_n585), .A3(new_n381), .A4(new_n328), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n329), .A2(G303), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n484), .A2(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n379), .A2(new_n381), .A3(new_n328), .A4(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n587), .C1(new_n589), .C2(KEYINPUT85), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n258), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n482), .A2(G270), .A3(new_n271), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n479), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n584), .A2(new_n596), .A3(G169), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n584), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(new_n595), .A3(G190), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n594), .A2(new_n479), .A3(G179), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n549), .A2(new_n605), .A3(new_n379), .A4(new_n588), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n591), .A3(new_n587), .A4(new_n586), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n607), .B2(new_n258), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n584), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n584), .A2(new_n596), .A3(KEYINPUT21), .A4(G169), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n599), .A2(new_n603), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n483), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n484), .A2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G250), .B2(G1698), .ZN(new_n614));
  INV_X1    g0414(.A(G294), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n382), .A2(new_n614), .B1(new_n325), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n612), .A2(G264), .B1(new_n616), .B2(new_n258), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n479), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n348), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n373), .A3(new_n479), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n519), .A2(G20), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT23), .B1(new_n222), .B2(G20), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT22), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n207), .A2(G87), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n329), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n385), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(KEYINPUT87), .C1(new_n543), .C2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n549), .A2(new_n207), .A3(new_n379), .A4(new_n631), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT87), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n627), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT24), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n630), .B1(new_n543), .B2(new_n632), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT24), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(new_n627), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n283), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT25), .B1(new_n318), .B2(new_n222), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n561), .A2(G107), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n622), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n642), .B2(new_n627), .ZN(new_n652));
  INV_X1    g0452(.A(new_n627), .ZN(new_n653));
  AOI211_X1 g0453(.A(KEYINPUT24), .B(new_n653), .C1(new_n641), .C2(new_n633), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n282), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n618), .A2(new_n436), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(G190), .B2(new_n618), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n649), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n567), .A2(new_n611), .A3(new_n651), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n459), .A2(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n350), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n430), .B(KEYINPUT18), .ZN(new_n662));
  OAI221_X1 g0462(.A(new_n454), .B1(new_n456), .B2(new_n453), .C1(new_n448), .C2(new_n449), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n280), .A2(new_n306), .ZN(new_n664));
  INV_X1    g0464(.A(new_n376), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n663), .A2(new_n303), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n440), .A2(new_n442), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n445), .B1(new_n667), .B2(KEYINPUT17), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n662), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n661), .B1(new_n670), .B2(new_n347), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n566), .B2(new_n504), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n527), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n522), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n563), .B(new_n564), .C1(new_n677), .C2(G169), .ZN(new_n678));
  INV_X1    g0478(.A(new_n504), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n546), .B(new_n556), .C1(new_n677), .C2(new_n436), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n672), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT90), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n672), .A2(new_n685), .A3(new_n682), .A4(new_n678), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n681), .A2(new_n678), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n504), .A2(new_n514), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n658), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n621), .B1(new_n655), .B2(new_n649), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n599), .A2(new_n609), .A3(new_n610), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n687), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n599), .A2(new_n609), .A3(new_n610), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n651), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n681), .A2(new_n678), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n515), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT89), .A4(new_n658), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n684), .A2(new_n686), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n671), .B1(new_n459), .B2(new_n700), .ZN(G369));
  NAND2_X1  g0501(.A1(new_n295), .A2(new_n207), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(G213), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n601), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n599), .A2(new_n603), .A3(new_n609), .A4(new_n610), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n651), .A2(new_n658), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n708), .B1(new_n655), .B2(new_n649), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(new_n651), .B2(new_n708), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n691), .A2(new_n708), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n651), .A2(new_n658), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n695), .A2(new_n707), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n719), .A3(new_n722), .ZN(G399));
  NAND2_X1  g0523(.A1(new_n210), .A2(new_n252), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n537), .A2(new_n385), .A3(new_n569), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n214), .B2(new_n724), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  INV_X1    g0530(.A(new_n678), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n566), .A2(new_n504), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n680), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n697), .B2(new_n504), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n734), .C1(new_n693), .C2(new_n690), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n730), .B1(new_n735), .B2(new_n708), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n684), .A2(new_n686), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n694), .A2(new_n699), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n707), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n736), .B1(new_n739), .B2(new_n730), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT91), .ZN(new_n741));
  AND4_X1   g0541(.A1(G244), .A2(new_n379), .A3(new_n381), .A4(new_n328), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G1698), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n550), .A3(new_n519), .A4(new_n552), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n527), .B1(new_n744), .B2(new_n258), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n608), .A3(new_n617), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n503), .A2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n745), .A2(new_n503), .A3(new_n608), .A4(new_n617), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n554), .A2(new_n617), .A3(new_n555), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n750), .B(new_n485), .C1(new_n471), .C2(new_n258), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT91), .A4(new_n608), .ZN(new_n754));
  INV_X1    g0554(.A(new_n503), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n554), .A2(new_n674), .A3(new_n675), .ZN(new_n756));
  AOI21_X1  g0556(.A(G179), .B1(new_n617), .B2(new_n479), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n755), .A2(new_n756), .A3(new_n596), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n748), .A2(new_n751), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n707), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n504), .A2(new_n514), .A3(new_n557), .A4(new_n565), .ZN(new_n765));
  NOR4_X1   g0565(.A1(new_n715), .A2(new_n711), .A3(new_n765), .A4(new_n707), .ZN(new_n766));
  OAI21_X1  g0566(.A(G330), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n762), .B(new_n763), .C1(new_n659), .C2(new_n707), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT92), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n770), .A3(G330), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n740), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n729), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n712), .A2(G330), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n294), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n206), .B1(new_n777), .B2(G45), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n776), .B(new_n714), .C1(new_n724), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n724), .ZN(new_n780));
  INV_X1    g0580(.A(new_n778), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n210), .A2(new_n261), .ZN(new_n783));
  INV_X1    g0583(.A(G355), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n784), .B1(G116), .B2(new_n210), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n243), .A2(G45), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n210), .A2(new_n382), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n253), .B2(new_n215), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(G20), .B1(KEYINPUT93), .B2(G169), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(KEYINPUT93), .A2(G169), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n216), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n782), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n207), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n615), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n207), .A2(new_n373), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(KEYINPUT33), .A2(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(KEYINPUT33), .A2(G317), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n804), .A2(new_n337), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n802), .B(new_n809), .C1(G326), .C2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n803), .A2(G190), .A3(new_n436), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n261), .B1(new_n813), .B2(G322), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G190), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n207), .A2(G179), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G311), .A2(new_n817), .B1(new_n820), .B2(G329), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n818), .A2(G190), .A3(G200), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(KEYINPUT95), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n818), .A2(new_n337), .A3(G200), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT96), .Z(new_n828));
  AOI22_X1  g0628(.A1(new_n826), .A2(G303), .B1(new_n828), .B2(G283), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n811), .A2(new_n814), .A3(new_n821), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n801), .A2(new_n489), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n261), .B1(new_n816), .B2(new_n220), .C1(new_n407), .C2(new_n812), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT32), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n819), .A2(new_n417), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n810), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(new_n202), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G68), .B2(new_n805), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n828), .A2(G107), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n826), .A2(G87), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n835), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n799), .B1(new_n842), .B2(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n796), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n712), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n779), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  NAND2_X1  g0648(.A1(new_n372), .A2(new_n707), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n369), .A2(new_n370), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n359), .B1(new_n337), .B2(new_n358), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n376), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT100), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT100), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n371), .A2(new_n854), .A3(new_n376), .A4(new_n849), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n739), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n853), .B(new_n855), .C1(new_n376), .C2(new_n708), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n739), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n782), .B1(new_n859), .B2(new_n772), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n772), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n793), .A2(new_n794), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n782), .B1(new_n863), .B2(G77), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT98), .Z(new_n865));
  AOI22_X1  g0665(.A1(new_n813), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n836), .B2(new_n867), .C1(new_n868), .C2(new_n806), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT34), .Z(new_n870));
  NAND2_X1  g0670(.A1(new_n826), .A2(G50), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n828), .A2(G68), .ZN(new_n872));
  INV_X1    g0672(.A(new_n801), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(G58), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n382), .B1(new_n820), .B2(G132), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n871), .A2(new_n872), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n810), .A2(G303), .B1(new_n817), .B2(G116), .ZN(new_n877));
  INV_X1    g0677(.A(G283), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n806), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n826), .A2(G107), .ZN(new_n881));
  INV_X1    g0681(.A(new_n831), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n828), .A2(G87), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n329), .B1(new_n812), .B2(new_n615), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(G311), .B2(new_n820), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n870), .A2(new_n876), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n865), .B1(new_n887), .B2(new_n793), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n858), .B2(new_n795), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n861), .A2(new_n889), .ZN(G384));
  NAND2_X1  g0690(.A1(new_n303), .A2(new_n707), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n309), .B2(new_n663), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n664), .A2(new_n891), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n458), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n376), .A2(new_n707), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n857), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n415), .A2(new_n282), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n419), .B1(new_n405), .B2(new_n403), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(KEYINPUT16), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n427), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n705), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n668), .B2(new_n662), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n396), .A2(new_n400), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n906), .B1(new_n910), .B2(new_n907), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n440), .A3(new_n442), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n440), .A2(new_n442), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n705), .B(KEYINPUT101), .Z(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n424), .B2(new_n427), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n430), .A2(KEYINPUT37), .A3(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(KEYINPUT37), .A2(new_n912), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n902), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(KEYINPUT38), .C1(new_n446), .C2(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n901), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT102), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n430), .B2(new_n444), .ZN(new_n927));
  OAI211_X1 g0727(.A(KEYINPUT102), .B(new_n439), .C1(new_n401), .C2(new_n428), .ZN(new_n928));
  INV_X1    g0728(.A(new_n915), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n920), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n668), .A2(new_n662), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n915), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n909), .A2(new_n917), .A3(new_n902), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n925), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n458), .A2(new_n707), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n918), .A2(new_n922), .A3(KEYINPUT39), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n433), .A2(new_n914), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n924), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n740), .A2(new_n459), .ZN(new_n943));
  INV_X1    g0743(.A(new_n671), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n942), .B(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G330), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n897), .A2(new_n769), .A3(new_n858), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n923), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n897), .A2(new_n769), .A3(new_n858), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n950), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n930), .A2(KEYINPUT37), .B1(new_n913), .B2(new_n916), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n929), .B1(new_n668), .B2(new_n662), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n902), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n922), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n949), .A2(new_n950), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n720), .A2(new_n611), .A3(new_n567), .A4(new_n708), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT31), .B1(new_n759), .B2(new_n707), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n459), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n947), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n957), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n946), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT103), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT103), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n946), .A2(new_n964), .B1(new_n206), .B2(new_n777), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(G116), .A3(new_n217), .A4(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT36), .Z(new_n973));
  OR3_X1    g0773(.A1(new_n214), .A2(new_n220), .A3(new_n408), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n202), .A2(G68), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n206), .B(G13), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n969), .A2(new_n973), .A3(new_n976), .ZN(G367));
  INV_X1    g0777(.A(new_n361), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n797), .B1(new_n238), .B2(new_n787), .C1(new_n210), .C2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G107), .A2(new_n873), .B1(new_n810), .B2(G311), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n489), .B2(new_n827), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n813), .A2(G303), .B1(new_n820), .B2(G317), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n878), .B2(new_n816), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n382), .B1(new_n806), .B2(new_n615), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n825), .B2(new_n569), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n826), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT110), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n825), .A2(new_n407), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n805), .A2(G159), .B1(new_n810), .B2(G143), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n329), .B1(new_n820), .B2(G137), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n813), .A2(G150), .B1(new_n817), .B2(G50), .ZN(new_n994));
  INV_X1    g0794(.A(new_n827), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n873), .A2(G68), .B1(new_n995), .B2(G77), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT47), .Z(new_n999));
  INV_X1    g0799(.A(new_n793), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n782), .B(new_n979), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT111), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT111), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n546), .A2(new_n708), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n688), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n678), .B2(new_n1004), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1002), .B(new_n1003), .C1(new_n844), .C2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n689), .B1(new_n513), .B2(new_n708), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n679), .A2(new_n707), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n722), .A2(new_n719), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT107), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT107), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1010), .B1(new_n722), .B2(new_n719), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT44), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n718), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT108), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT108), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n722), .B1(new_n717), .B2(new_n721), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(new_n713), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n774), .A2(KEYINPUT109), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n772), .A3(new_n740), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n774), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n724), .B(KEYINPUT41), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n781), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1010), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n722), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT42), .ZN(new_n1042));
  XOR2_X1   g0842(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n1043));
  NOR2_X1   g0843(.A1(new_n1006), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n504), .B1(new_n1008), .B2(new_n651), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n708), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT105), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1021), .A2(new_n1010), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT106), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1044), .B1(KEYINPUT43), .B2(new_n1006), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1050), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1007), .B1(new_n1039), .B2(new_n1057), .ZN(G387));
  AND2_X1   g0858(.A1(new_n1032), .A2(new_n780), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n774), .B2(new_n1030), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n717), .A2(new_n844), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n783), .A2(new_n726), .B1(G107), .B2(new_n210), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n235), .A2(new_n253), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n310), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI211_X1 g0865(.A(G45), .B(new_n725), .C1(G68), .C2(G77), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n787), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1062), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n782), .B1(new_n1068), .B2(new_n798), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n361), .A2(new_n873), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n813), .A2(G50), .B1(new_n820), .B2(G150), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n289), .C2(new_n816), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n534), .B1(new_n836), .B2(new_n417), .C1(new_n310), .C2(new_n806), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n826), .A2(G77), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n828), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1074), .B(new_n1075), .C1(new_n489), .C2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n813), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n805), .A2(G311), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n810), .A2(G322), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n826), .A2(G294), .B1(G283), .B2(new_n873), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT112), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT49), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n534), .B1(G326), .B2(new_n820), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(new_n569), .C2(new_n827), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1087), .A2(KEYINPUT49), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1077), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1069), .B1(new_n1092), .B2(new_n793), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1030), .A2(new_n781), .B1(new_n1061), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1060), .A2(new_n1094), .ZN(G393));
  NAND2_X1  g0895(.A1(new_n1026), .A2(new_n1022), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n778), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1040), .A2(new_n796), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n246), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n797), .B1(new_n489), .B2(new_n210), .C1(new_n1099), .C2(new_n787), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n782), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n311), .A2(new_n817), .B1(new_n820), .B2(G143), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G77), .A2(new_n873), .B1(new_n805), .B2(G50), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n883), .A2(new_n534), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n810), .B1(new_n813), .B2(G159), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n826), .A2(G68), .B1(new_n1105), .B2(KEYINPUT51), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(KEYINPUT51), .B2(new_n1105), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G317), .A2(new_n810), .B1(new_n813), .B2(G311), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n826), .A2(G283), .B1(new_n1108), .B2(KEYINPUT52), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(KEYINPUT52), .B2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n329), .B1(new_n816), .B2(new_n615), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G322), .B2(new_n820), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G116), .A2(new_n873), .B1(new_n805), .B2(G303), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n839), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1104), .A2(new_n1107), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1101), .B1(new_n1115), .B2(new_n793), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1098), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1035), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1118), .A2(new_n1025), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n724), .B1(new_n1096), .B2(new_n1032), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(G390));
  INV_X1    g0922(.A(KEYINPUT113), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n856), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n700), .A2(new_n707), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n897), .B1(new_n1125), .B2(new_n899), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n938), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1126), .A2(new_n1127), .B1(new_n937), .B2(new_n939), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n938), .B1(new_n955), .B2(new_n922), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n732), .A2(new_n680), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n678), .A3(new_n734), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n690), .A2(new_n693), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n708), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n900), .B1(new_n1133), .B2(new_n1124), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n897), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n768), .A2(new_n771), .A3(new_n858), .A4(new_n897), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1123), .B1(new_n1128), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n937), .A2(new_n939), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n901), .B2(new_n938), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT113), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1136), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n947), .B1(new_n961), .B2(new_n958), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n897), .A2(new_n1145), .A3(new_n858), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1139), .A2(new_n1143), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n781), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1140), .A2(new_n794), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n782), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n862), .B2(new_n310), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  AOI22_X1  g0952(.A1(new_n873), .A2(G159), .B1(new_n817), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n867), .B2(new_n806), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT114), .Z(new_n1155));
  OR3_X1    g0955(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n868), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT53), .B1(new_n825), .B2(new_n868), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n261), .B1(new_n819), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G132), .B2(new_n813), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n810), .A2(G128), .B1(new_n995), .B2(G50), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1155), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G77), .A2(new_n873), .B1(new_n810), .B2(G283), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n222), .B2(new_n806), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n329), .B1(new_n812), .B2(new_n569), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n816), .A2(new_n489), .B1(new_n819), .B2(new_n615), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n840), .A2(new_n872), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1149), .B(new_n1151), .C1(new_n1000), .C2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1145), .A2(new_n446), .A3(new_n458), .A4(new_n378), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n671), .B(new_n1172), .C1(new_n740), .C2(new_n459), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1125), .A2(new_n899), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(KEYINPUT92), .B(new_n947), .C1(new_n961), .C2(new_n958), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n770), .B1(new_n769), .B2(G330), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n897), .B1(new_n1178), .B2(new_n858), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1179), .B2(new_n1146), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1145), .A2(new_n858), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1134), .B1(new_n898), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1137), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1173), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n780), .B1(new_n1147), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1136), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1146), .B1(new_n1128), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1128), .A2(new_n1123), .A3(new_n1138), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT113), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1184), .B(new_n1187), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1148), .B(new_n1171), .C1(new_n1185), .C2(new_n1191), .ZN(G378));
  INV_X1    g0992(.A(KEYINPUT120), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1173), .B1(new_n1147), .B2(new_n1184), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n705), .B1(new_n315), .B2(new_n319), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT55), .Z(new_n1197));
  XNOR2_X1  g0997(.A(new_n351), .B(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1199));
  XOR2_X1   g0999(.A(new_n1198), .B(new_n1199), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT119), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n957), .A2(G330), .A3(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n918), .A2(new_n922), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n950), .B1(new_n1203), .B2(new_n951), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n948), .A2(KEYINPUT40), .A3(new_n956), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(G330), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1200), .A2(KEYINPUT119), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n942), .A2(new_n1202), .A3(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n901), .A2(new_n923), .B1(new_n433), .B2(new_n914), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1202), .A2(new_n1208), .B1(new_n940), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1194), .B1(new_n1195), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1173), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1190), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n940), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1201), .B1(new_n957), .B2(G330), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n942), .A2(new_n1202), .A3(new_n1208), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1194), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n724), .B1(new_n1215), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1213), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n781), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1200), .A2(new_n794), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n782), .B1(new_n863), .B2(G50), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n805), .A2(G132), .ZN(new_n1227));
  INV_X1    g1027(.A(G128), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n812), .C1(new_n867), .C2(new_n816), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n836), .A2(new_n1158), .B1(new_n868), .B2(new_n801), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT116), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(new_n826), .C2(new_n1152), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT59), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n820), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n325), .A3(new_n252), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G159), .B2(new_n995), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n827), .A2(new_n407), .B1(new_n819), .B2(new_n878), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n382), .A2(new_n252), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1075), .A2(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT115), .Z(new_n1246));
  OAI22_X1  g1046(.A1(new_n801), .A2(new_n289), .B1(new_n812), .B2(new_n222), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n806), .A2(new_n489), .B1(new_n836), .B2(new_n569), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n361), .C2(new_n817), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1240), .A2(new_n1241), .B1(KEYINPUT58), .B2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1243), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(KEYINPUT58), .C2(new_n1250), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1226), .B1(new_n1253), .B2(new_n793), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1225), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1224), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1193), .B1(new_n1223), .B2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(KEYINPUT120), .B(new_n1256), .C1(new_n1213), .C2(new_n1222), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(G375));
  INV_X1    g1060(.A(new_n1184), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n768), .A2(new_n771), .A3(new_n858), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1146), .B1(new_n1262), .B2(new_n898), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1173), .B(new_n1183), .C1(new_n1263), .C2(new_n1174), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1038), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1183), .B1(new_n1263), .B2(new_n1174), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n781), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n863), .A2(G68), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1076), .A2(new_n220), .B1(new_n825), .B2(new_n489), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n805), .A2(G116), .B1(new_n810), .B2(G294), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n261), .B1(new_n813), .B2(G283), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G107), .A2(new_n817), .B1(new_n820), .B2(G303), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(new_n1070), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n825), .A2(new_n417), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n816), .A2(new_n868), .B1(new_n819), .B2(new_n1228), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G137), .B2(new_n813), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G50), .A2(new_n873), .B1(new_n810), .B2(G132), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n805), .A2(new_n1152), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n382), .B1(new_n995), .B2(G58), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1269), .A2(new_n1273), .B1(new_n1274), .B2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1150), .B(new_n1268), .C1(new_n1281), .C2(new_n793), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n897), .B2(new_n795), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1267), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1265), .A2(new_n1285), .ZN(G381));
  OAI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n780), .B1(new_n1195), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1257), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT120), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1223), .A2(new_n1193), .A3(new_n1257), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G378), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1037), .B1(new_n1119), .B2(new_n774), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1056), .B1(new_n1295), .B2(new_n781), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1060), .A2(new_n847), .A3(new_n1094), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G390), .A2(G381), .A3(new_n1297), .A4(G384), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1294), .A2(new_n1007), .A3(new_n1296), .A4(new_n1298), .ZN(G407));
  OAI21_X1  g1099(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1171), .B1(new_n1300), .B2(new_n778), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n724), .B1(new_n1300), .B2(new_n1261), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1190), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G407), .B(G213), .C1(G343), .C2(new_n1304), .ZN(G409));
  INV_X1    g1105(.A(new_n1297), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n847), .B1(new_n1060), .B2(new_n1094), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G390), .B(new_n1007), .C1(new_n1039), .C2(new_n1057), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1296), .B2(new_n1007), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G387), .A2(new_n1121), .A3(new_n1117), .ZN(new_n1313));
  OR3_X1    g1113(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1308), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1315), .A3(new_n1309), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n706), .A2(G213), .ZN(new_n1318));
  INV_X1    g1118(.A(G2897), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(KEYINPUT124), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(KEYINPUT124), .B2(new_n1319), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n724), .B1(new_n1266), .B2(new_n1214), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1264), .A2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n1173), .A4(new_n1183), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1322), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT121), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1322), .A2(new_n1324), .A3(new_n1325), .A4(KEYINPUT121), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1285), .ZN(new_n1331));
  INV_X1    g1131(.A(G384), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(G384), .A3(new_n1285), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT122), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G384), .B1(new_n1330), .B2(new_n1285), .ZN(new_n1336));
  AOI211_X1 g1136(.A(new_n1332), .B(new_n1284), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT122), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1321), .B1(new_n1335), .B2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1318), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(G2897), .A3(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1340), .A2(KEYINPUT125), .A3(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT125), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1321), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1333), .A2(KEYINPUT122), .A3(new_n1334), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1338), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1347), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1341), .A2(new_n1319), .A3(new_n1318), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1346), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  OAI211_X1 g1152(.A(G378), .B(new_n1257), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1195), .A2(new_n1212), .A3(new_n1037), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1303), .B1(new_n1354), .B2(new_n1256), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1343), .B1(new_n1353), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1345), .A2(new_n1352), .A3(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT61), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1356), .A2(new_n1360), .A3(KEYINPUT62), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT62), .B1(new_n1356), .B2(new_n1360), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1359), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1317), .B1(new_n1358), .B2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1356), .A2(new_n1360), .A3(KEYINPUT63), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1365), .A2(new_n1366), .A3(new_n1359), .ZN(new_n1367));
  AOI21_X1  g1167(.A(KEYINPUT63), .B1(new_n1356), .B2(new_n1360), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(new_n1356), .B(KEYINPUT123), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1370), .A2(new_n1352), .A3(new_n1345), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1364), .A2(new_n1372), .ZN(G405));
  NAND2_X1  g1173(.A1(new_n1291), .A2(G378), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1342), .B1(new_n1294), .B2(new_n1375), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1304), .A2(new_n1360), .A3(new_n1374), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1376), .A2(new_n1377), .A3(new_n1317), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT127), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1381), .A2(new_n1366), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1376), .A2(new_n1377), .A3(new_n1317), .A4(KEYINPUT127), .ZN(new_n1383));
  AND3_X1   g1183(.A1(new_n1380), .A2(new_n1382), .A3(new_n1383), .ZN(G402));
endmodule


