

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X2 U551 ( .A(KEYINPUT68), .B(n522), .Z(n897) );
  XOR2_X2 U552 ( .A(KEYINPUT17), .B(n521), .Z(n892) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n656) );
  INV_X1 U554 ( .A(n643), .ZN(n638) );
  XNOR2_X1 U555 ( .A(n635), .B(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U556 ( .A(n637), .B(n636), .ZN(n642) );
  XNOR2_X1 U557 ( .A(n657), .B(n656), .ZN(n666) );
  NOR2_X2 U558 ( .A1(n518), .A2(G2105), .ZN(n893) );
  INV_X1 U559 ( .A(KEYINPUT40), .ZN(n758) );
  NOR2_X1 U560 ( .A1(G651), .A2(n556), .ZN(n791) );
  XNOR2_X1 U561 ( .A(n758), .B(KEYINPUT105), .ZN(n759) );
  XNOR2_X1 U562 ( .A(n587), .B(KEYINPUT65), .ZN(n589) );
  XOR2_X1 U563 ( .A(G2104), .B(KEYINPUT66), .Z(n518) );
  NAND2_X1 U564 ( .A1(G102), .A2(n893), .ZN(n520) );
  AND2_X1 U565 ( .A1(G2105), .A2(n518), .ZN(n896) );
  NAND2_X1 U566 ( .A1(G126), .A2(n896), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NAND2_X1 U569 ( .A1(G138), .A2(n892), .ZN(n524) );
  NAND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  NAND2_X1 U571 ( .A1(G114), .A2(n897), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U573 ( .A1(n526), .A2(n525), .ZN(G164) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n556) );
  NAND2_X1 U575 ( .A1(n791), .A2(G52), .ZN(n529) );
  XOR2_X1 U576 ( .A(G651), .B(KEYINPUT72), .Z(n530) );
  NOR2_X1 U577 ( .A1(G543), .A2(n530), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n527), .Z(n792) );
  NAND2_X1 U579 ( .A1(G64), .A2(n792), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n795) );
  NAND2_X1 U582 ( .A1(n795), .A2(G90), .ZN(n532) );
  NOR2_X1 U583 ( .A1(n556), .A2(n530), .ZN(n796) );
  NAND2_X1 U584 ( .A1(G77), .A2(n796), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(n533), .Z(n534) );
  NOR2_X1 U587 ( .A1(n535), .A2(n534), .ZN(G171) );
  NAND2_X1 U588 ( .A1(n795), .A2(G88), .ZN(n537) );
  NAND2_X1 U589 ( .A1(G75), .A2(n796), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n792), .A2(G62), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT86), .B(n538), .Z(n539) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n791), .A2(G50), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(G303) );
  NAND2_X1 U596 ( .A1(n791), .A2(G51), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G63), .A2(n792), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT6), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n546), .B(KEYINPUT79), .ZN(n553) );
  XNOR2_X1 U601 ( .A(KEYINPUT78), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n795), .A2(G89), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G76), .A2(n796), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U608 ( .A(KEYINPUT7), .B(n554), .ZN(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U610 ( .A1(G74), .A2(G651), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n555), .B(KEYINPUT84), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G49), .A2(n791), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G87), .A2(n556), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U615 ( .A1(n792), .A2(n559), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(G288) );
  NAND2_X1 U617 ( .A1(G61), .A2(n792), .ZN(n568) );
  NAND2_X1 U618 ( .A1(G86), .A2(n795), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G48), .A2(n791), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n796), .A2(G73), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT2), .B(n564), .Z(n565) );
  NOR2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT85), .B(n569), .Z(G305) );
  NAND2_X1 U626 ( .A1(n795), .A2(G85), .ZN(n571) );
  NAND2_X1 U627 ( .A1(G72), .A2(n796), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n791), .A2(G47), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G60), .A2(n792), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U632 ( .A1(n575), .A2(n574), .ZN(G290) );
  NAND2_X1 U633 ( .A1(n892), .A2(G137), .ZN(n576) );
  XNOR2_X1 U634 ( .A(n576), .B(KEYINPUT70), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G113), .A2(n897), .ZN(n577) );
  XOR2_X1 U636 ( .A(n577), .B(KEYINPUT69), .Z(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U638 ( .A(n580), .B(KEYINPUT71), .ZN(n586) );
  NAND2_X1 U639 ( .A1(n893), .A2(G101), .ZN(n581) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n581), .Z(n583) );
  NAND2_X1 U641 ( .A1(n896), .A2(G125), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U643 ( .A(n584), .B(KEYINPUT67), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n587) );
  BUF_X1 U645 ( .A(n589), .Z(G160) );
  NOR2_X1 U646 ( .A1(G164), .A2(G1384), .ZN(n692) );
  AND2_X1 U647 ( .A1(G40), .A2(n692), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U649 ( .A(n590), .B(KEYINPUT64), .ZN(n643) );
  NAND2_X1 U650 ( .A1(G2072), .A2(n638), .ZN(n591) );
  XNOR2_X1 U651 ( .A(n591), .B(KEYINPUT27), .ZN(n593) );
  INV_X1 U652 ( .A(G1956), .ZN(n943) );
  NOR2_X1 U653 ( .A1(n638), .A2(n943), .ZN(n592) );
  NOR2_X1 U654 ( .A1(n593), .A2(n592), .ZN(n601) );
  NAND2_X1 U655 ( .A1(n791), .A2(G53), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G65), .A2(n792), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n795), .A2(G91), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G78), .A2(n796), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U661 ( .A1(n599), .A2(n598), .ZN(n1004) );
  NOR2_X1 U662 ( .A1(n601), .A2(n1004), .ZN(n600) );
  XOR2_X1 U663 ( .A(n600), .B(KEYINPUT28), .Z(n634) );
  NAND2_X1 U664 ( .A1(n601), .A2(n1004), .ZN(n632) );
  NAND2_X1 U665 ( .A1(G54), .A2(n791), .ZN(n608) );
  NAND2_X1 U666 ( .A1(G79), .A2(n796), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G66), .A2(n792), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n795), .A2(G92), .ZN(n604) );
  XOR2_X1 U670 ( .A(KEYINPUT76), .B(n604), .Z(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U672 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U673 ( .A(n609), .B(KEYINPUT15), .ZN(n1010) );
  NAND2_X1 U674 ( .A1(n638), .A2(G1996), .ZN(n610) );
  XNOR2_X1 U675 ( .A(n610), .B(KEYINPUT26), .ZN(n623) );
  AND2_X1 U676 ( .A1(n643), .A2(G1341), .ZN(n621) );
  NAND2_X1 U677 ( .A1(G56), .A2(n792), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n611), .Z(n617) );
  NAND2_X1 U679 ( .A1(n795), .A2(G81), .ZN(n612) );
  XNOR2_X1 U680 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G68), .A2(n796), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U685 ( .A(n618), .B(KEYINPUT74), .ZN(n620) );
  NAND2_X1 U686 ( .A1(G43), .A2(n791), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n1018) );
  NOR2_X1 U688 ( .A1(n621), .A2(n1018), .ZN(n622) );
  AND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n628) );
  NOR2_X1 U690 ( .A1(n1010), .A2(n628), .ZN(n627) );
  NAND2_X1 U691 ( .A1(G2067), .A2(n638), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n643), .A2(G1348), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n630) );
  AND2_X1 U695 ( .A1(n628), .A2(n1010), .ZN(n629) );
  NOR2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U698 ( .A1(n634), .A2(n633), .ZN(n637) );
  INV_X1 U699 ( .A(KEYINPUT100), .ZN(n635) );
  XNOR2_X1 U700 ( .A(KEYINPUT25), .B(G2078), .ZN(n926) );
  NOR2_X1 U701 ( .A1(n643), .A2(n926), .ZN(n640) );
  INV_X1 U702 ( .A(G1961), .ZN(n941) );
  NOR2_X1 U703 ( .A1(n638), .A2(n941), .ZN(n639) );
  NOR2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n653) );
  NAND2_X1 U705 ( .A1(n653), .A2(G171), .ZN(n641) );
  NAND2_X1 U706 ( .A1(n642), .A2(n641), .ZN(n665) );
  INV_X1 U707 ( .A(G8), .ZN(n648) );
  NOR2_X1 U708 ( .A1(n643), .A2(G2090), .ZN(n645) );
  NAND2_X1 U709 ( .A1(n643), .A2(G8), .ZN(n734) );
  NOR2_X1 U710 ( .A1(G1971), .A2(n734), .ZN(n644) );
  NOR2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n646), .A2(G303), .ZN(n647) );
  OR2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n659) );
  AND2_X1 U714 ( .A1(n665), .A2(n659), .ZN(n658) );
  NOR2_X1 U715 ( .A1(n734), .A2(G1966), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n649), .B(KEYINPUT99), .ZN(n669) );
  NOR2_X1 U717 ( .A1(n643), .A2(G2084), .ZN(n667) );
  NOR2_X1 U718 ( .A1(n648), .A2(n667), .ZN(n650) );
  AND2_X1 U719 ( .A1(n669), .A2(n650), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT30), .B(n651), .Z(n652) );
  NOR2_X1 U721 ( .A1(G168), .A2(n652), .ZN(n655) );
  NOR2_X1 U722 ( .A1(G171), .A2(n653), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n666), .ZN(n663) );
  INV_X1 U725 ( .A(n659), .ZN(n661) );
  AND2_X1 U726 ( .A1(G286), .A2(G8), .ZN(n660) );
  OR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U729 ( .A(n664), .B(KEYINPUT32), .ZN(n725) );
  NAND2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n671) );
  NAND2_X1 U731 ( .A1(G8), .A2(n667), .ZN(n668) );
  AND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n723) );
  NAND2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n1016) );
  AND2_X1 U735 ( .A1(n723), .A2(n1016), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n725), .A2(n672), .ZN(n716) );
  INV_X1 U737 ( .A(n1016), .ZN(n674) );
  NOR2_X1 U738 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n1007) );
  NOR2_X1 U740 ( .A1(n1013), .A2(n1007), .ZN(n673) );
  OR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n714) );
  NAND2_X1 U742 ( .A1(n1013), .A2(KEYINPUT33), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n675), .A2(n734), .ZN(n677) );
  XOR2_X1 U744 ( .A(G1981), .B(G305), .Z(n1028) );
  INV_X1 U745 ( .A(n1028), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n712) );
  NAND2_X1 U747 ( .A1(G140), .A2(n892), .ZN(n679) );
  NAND2_X1 U748 ( .A1(G104), .A2(n893), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(KEYINPUT93), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT34), .ZN(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n685) );
  NAND2_X1 U753 ( .A1(G128), .A2(n896), .ZN(n683) );
  NAND2_X1 U754 ( .A1(G116), .A2(n897), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U758 ( .A(KEYINPUT36), .B(n688), .Z(n875) );
  XNOR2_X1 U759 ( .A(G2067), .B(KEYINPUT37), .ZN(n689) );
  XNOR2_X1 U760 ( .A(n689), .B(KEYINPUT92), .ZN(n752) );
  NOR2_X1 U761 ( .A1(n875), .A2(n752), .ZN(n690) );
  XNOR2_X1 U762 ( .A(n690), .B(KEYINPUT95), .ZN(n980) );
  XOR2_X1 U763 ( .A(G1986), .B(G290), .Z(n1009) );
  NAND2_X1 U764 ( .A1(n980), .A2(n1009), .ZN(n693) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n754) );
  AND2_X1 U767 ( .A1(n693), .A2(n754), .ZN(n711) );
  NAND2_X1 U768 ( .A1(G141), .A2(n892), .ZN(n695) );
  NAND2_X1 U769 ( .A1(G129), .A2(n896), .ZN(n694) );
  NAND2_X1 U770 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n893), .A2(G105), .ZN(n696) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(n696), .Z(n697) );
  NOR2_X1 U773 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U774 ( .A1(G117), .A2(n897), .ZN(n699) );
  NAND2_X1 U775 ( .A1(n700), .A2(n699), .ZN(n874) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n874), .ZN(n701) );
  XNOR2_X1 U777 ( .A(n701), .B(KEYINPUT97), .ZN(n709) );
  XOR2_X1 U778 ( .A(KEYINPUT96), .B(G1991), .Z(n922) );
  NAND2_X1 U779 ( .A1(G131), .A2(n892), .ZN(n703) );
  NAND2_X1 U780 ( .A1(G119), .A2(n896), .ZN(n702) );
  NAND2_X1 U781 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U782 ( .A1(G95), .A2(n893), .ZN(n705) );
  NAND2_X1 U783 ( .A1(G107), .A2(n897), .ZN(n704) );
  NAND2_X1 U784 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n903) );
  NOR2_X1 U786 ( .A1(n922), .A2(n903), .ZN(n708) );
  NOR2_X1 U787 ( .A1(n709), .A2(n708), .ZN(n987) );
  INV_X1 U788 ( .A(n754), .ZN(n710) );
  NOR2_X1 U789 ( .A1(n987), .A2(n710), .ZN(n746) );
  NOR2_X1 U790 ( .A1(n711), .A2(n746), .ZN(n737) );
  AND2_X1 U791 ( .A1(n712), .A2(n737), .ZN(n717) );
  AND2_X1 U792 ( .A1(n717), .A2(KEYINPUT33), .ZN(n720) );
  INV_X1 U793 ( .A(n720), .ZN(n713) );
  AND2_X1 U794 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U795 ( .A1(n716), .A2(n715), .ZN(n722) );
  INV_X1 U796 ( .A(n717), .ZN(n718) );
  NOR2_X1 U797 ( .A1(n734), .A2(n718), .ZN(n719) );
  OR2_X1 U798 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n722), .A2(n721), .ZN(n741) );
  AND2_X1 U800 ( .A1(n734), .A2(n737), .ZN(n726) );
  AND2_X1 U801 ( .A1(n723), .A2(n726), .ZN(n724) );
  NAND2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n731) );
  INV_X1 U803 ( .A(n726), .ZN(n729) );
  NOR2_X1 U804 ( .A1(G2090), .A2(G303), .ZN(n727) );
  NAND2_X1 U805 ( .A1(G8), .A2(n727), .ZN(n728) );
  OR2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n739) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n732) );
  XOR2_X1 U809 ( .A(n732), .B(KEYINPUT98), .Z(n733) );
  XNOR2_X1 U810 ( .A(KEYINPUT24), .B(n733), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  INV_X1 U815 ( .A(KEYINPUT102), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n743), .B(n742), .ZN(n757) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n874), .ZN(n978) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n744) );
  AND2_X1 U819 ( .A1(n922), .A2(n903), .ZN(n989) );
  NOR2_X1 U820 ( .A1(n744), .A2(n989), .ZN(n745) );
  NOR2_X1 U821 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U822 ( .A(KEYINPUT103), .B(n747), .Z(n748) );
  NOR2_X1 U823 ( .A1(n978), .A2(n748), .ZN(n749) );
  XNOR2_X1 U824 ( .A(n749), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n750), .A2(n980), .ZN(n751) );
  XNOR2_X1 U826 ( .A(n751), .B(KEYINPUT104), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n752), .A2(n875), .ZN(n990) );
  NAND2_X1 U828 ( .A1(n753), .A2(n990), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n760) );
  XNOR2_X1 U831 ( .A(n760), .B(n759), .ZN(G329) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G123), .A2(n896), .ZN(n761) );
  XNOR2_X1 U834 ( .A(n761), .B(KEYINPUT18), .ZN(n768) );
  NAND2_X1 U835 ( .A1(G135), .A2(n892), .ZN(n763) );
  NAND2_X1 U836 ( .A1(G111), .A2(n897), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U838 ( .A1(G99), .A2(n893), .ZN(n764) );
  XNOR2_X1 U839 ( .A(KEYINPUT83), .B(n764), .ZN(n765) );
  NOR2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n986) );
  XNOR2_X1 U842 ( .A(G2096), .B(n986), .ZN(n769) );
  OR2_X1 U843 ( .A1(G2100), .A2(n769), .ZN(G156) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U846 ( .A(n770), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U847 ( .A(G223), .ZN(n839) );
  NAND2_X1 U848 ( .A1(n839), .A2(G567), .ZN(n771) );
  XNOR2_X1 U849 ( .A(n771), .B(KEYINPUT11), .ZN(n772) );
  XNOR2_X1 U850 ( .A(KEYINPUT73), .B(n772), .ZN(G234) );
  INV_X1 U851 ( .A(G860), .ZN(n790) );
  OR2_X1 U852 ( .A1(n1018), .A2(n790), .ZN(G153) );
  INV_X1 U853 ( .A(G868), .ZN(n783) );
  NOR2_X1 U854 ( .A1(n783), .A2(G171), .ZN(n773) );
  XNOR2_X1 U855 ( .A(n773), .B(KEYINPUT75), .ZN(n775) );
  INV_X1 U856 ( .A(n1010), .ZN(n784) );
  NAND2_X1 U857 ( .A1(n783), .A2(n784), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U859 ( .A(KEYINPUT77), .B(n776), .Z(G284) );
  INV_X1 U860 ( .A(n1004), .ZN(G299) );
  NOR2_X1 U861 ( .A1(G868), .A2(G299), .ZN(n777) );
  XNOR2_X1 U862 ( .A(n777), .B(KEYINPUT80), .ZN(n779) );
  NOR2_X1 U863 ( .A1(n783), .A2(G286), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U865 ( .A1(G559), .A2(n790), .ZN(n780) );
  XOR2_X1 U866 ( .A(KEYINPUT81), .B(n780), .Z(n781) );
  NAND2_X1 U867 ( .A1(n781), .A2(n1010), .ZN(n782) );
  XNOR2_X1 U868 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U870 ( .A(KEYINPUT82), .B(n785), .Z(n786) );
  NOR2_X1 U871 ( .A1(G559), .A2(n786), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G868), .A2(n1018), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G559), .A2(n1010), .ZN(n789) );
  XOR2_X1 U875 ( .A(n1018), .B(n789), .Z(n808) );
  NAND2_X1 U876 ( .A1(n790), .A2(n808), .ZN(n801) );
  NAND2_X1 U877 ( .A1(n791), .A2(G55), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G67), .A2(n792), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U880 ( .A1(n795), .A2(G93), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G80), .A2(n796), .ZN(n797) );
  NAND2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n810) );
  XOR2_X1 U884 ( .A(n801), .B(n810), .Z(G145) );
  INV_X1 U885 ( .A(G303), .ZN(G166) );
  XOR2_X1 U886 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n802) );
  XNOR2_X1 U887 ( .A(G288), .B(n802), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n810), .B(n803), .ZN(n805) );
  XNOR2_X1 U889 ( .A(G290), .B(n1004), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U891 ( .A(n806), .B(G305), .Z(n807) );
  XNOR2_X1 U892 ( .A(G166), .B(n807), .ZN(n910) );
  XNOR2_X1 U893 ( .A(n808), .B(n910), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n809), .A2(G868), .ZN(n812) );
  OR2_X1 U895 ( .A1(G868), .A2(n810), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n814), .ZN(n816) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(KEYINPUT88), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U902 ( .A1(G2072), .A2(n817), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n819) );
  NAND2_X1 U905 ( .A1(G132), .A2(G82), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n819), .B(n818), .ZN(n820) );
  NOR2_X1 U907 ( .A1(n820), .A2(G218), .ZN(n821) );
  NAND2_X1 U908 ( .A1(G96), .A2(n821), .ZN(n845) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n845), .ZN(n825) );
  NAND2_X1 U910 ( .A1(G69), .A2(G120), .ZN(n822) );
  NOR2_X1 U911 ( .A1(G237), .A2(n822), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G108), .A2(n823), .ZN(n846) );
  NAND2_X1 U913 ( .A1(G567), .A2(n846), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U915 ( .A(KEYINPUT90), .B(n826), .ZN(n865) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n865), .A2(n827), .ZN(n844) );
  NAND2_X1 U918 ( .A1(G36), .A2(n844), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT91), .B(n828), .Z(G176) );
  XNOR2_X1 U920 ( .A(KEYINPUT106), .B(G2454), .ZN(n837) );
  XNOR2_X1 U921 ( .A(G2430), .B(G2435), .ZN(n835) );
  XOR2_X1 U922 ( .A(G2451), .B(G2427), .Z(n830) );
  XNOR2_X1 U923 ( .A(G2438), .B(G2446), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U925 ( .A(n831), .B(G2443), .Z(n833) );
  XNOR2_X1 U926 ( .A(G1348), .B(G1341), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n838), .A2(G14), .ZN(n915) );
  XNOR2_X1 U931 ( .A(KEYINPUT107), .B(n915), .ZN(G401) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n839), .ZN(G217) );
  INV_X1 U933 ( .A(G661), .ZN(n841) );
  NAND2_X1 U934 ( .A1(G2), .A2(G15), .ZN(n840) );
  NOR2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U936 ( .A(KEYINPUT108), .B(n842), .Z(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U940 ( .A(G132), .ZN(G219) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U947 ( .A(G1991), .B(KEYINPUT41), .ZN(n856) );
  XOR2_X1 U948 ( .A(G1971), .B(G1956), .Z(n848) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1986), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n850) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U953 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U954 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U955 ( .A(G2474), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n860) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(G227) );
  XNOR2_X1 U967 ( .A(KEYINPUT109), .B(n865), .ZN(G319) );
  NAND2_X1 U968 ( .A1(G100), .A2(n893), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G112), .A2(n897), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G124), .A2(n896), .ZN(n868) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n868), .Z(n869) );
  XNOR2_X1 U973 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G136), .A2(n892), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U977 ( .A(n875), .B(n874), .Z(n876) );
  XNOR2_X1 U978 ( .A(n986), .B(n876), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G130), .A2(n896), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G118), .A2(n897), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G142), .A2(n892), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G106), .A2(n893), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n881), .Z(n882) );
  NOR2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U988 ( .A(G164), .B(G162), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U990 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n889) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U992 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U993 ( .A(n891), .B(n890), .Z(n905) );
  NAND2_X1 U994 ( .A1(G139), .A2(n892), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n982) );
  XNOR2_X1 U1002 ( .A(n903), .B(n982), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(G160), .B(n906), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(n1018), .B(G286), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(G171), .B(n1010), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  XNOR2_X1 U1011 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n915), .A2(G319), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT114), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n917) );
  XOR2_X1 U1017 ( .A(KEYINPUT116), .B(n917), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1022 ( .A(n922), .B(G25), .Z(n924) );
  XNOR2_X1 U1023 ( .A(G2067), .B(G26), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G2072), .B(G33), .Z(n925) );
  NAND2_X1 U1026 ( .A1(G28), .A2(n925), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G1996), .B(G32), .Z(n928) );
  XNOR2_X1 U1028 ( .A(n926), .B(G27), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1030 ( .A(KEYINPUT117), .B(n929), .Z(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT53), .ZN(n937) );
  XOR2_X1 U1034 ( .A(G2084), .B(KEYINPUT54), .Z(n935) );
  XNOR2_X1 U1035 ( .A(G34), .B(n935), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n970) );
  NAND2_X1 U1039 ( .A1(KEYINPUT55), .A2(n970), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n940), .ZN(n976) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT122), .ZN(n968) );
  XNOR2_X1 U1042 ( .A(n941), .B(G5), .ZN(n964) );
  XOR2_X1 U1043 ( .A(G1966), .B(KEYINPUT124), .Z(n942) );
  XNOR2_X1 U1044 ( .A(G21), .B(n942), .ZN(n954) );
  XOR2_X1 U1045 ( .A(G1341), .B(G19), .Z(n945) );
  XNOR2_X1 U1046 ( .A(n943), .B(G20), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G1981), .B(G6), .Z(n949) );
  XOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT123), .Z(n946) );
  XNOR2_X1 U1050 ( .A(G4), .B(n946), .ZN(n947) );
  XNOR2_X1 U1051 ( .A(n947), .B(KEYINPUT59), .ZN(n948) );
  NAND2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1054 ( .A(n952), .B(KEYINPUT60), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n960) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n958) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n956) );
  XNOR2_X1 U1059 ( .A(G23), .B(G1976), .ZN(n955) );
  NOR2_X1 U1060 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1062 ( .A(n960), .B(n959), .Z(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(n965), .B(KEYINPUT61), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(n966), .B(KEYINPUT126), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(KEYINPUT127), .B(n969), .ZN(n974) );
  INV_X1 U1069 ( .A(n970), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(G29), .A2(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n1003) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n979), .Z(n981) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n997) );
  XOR2_X1 U1078 ( .A(G2072), .B(n982), .Z(n984) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT50), .B(n985), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1085 ( .A(G160), .B(G2084), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(n998), .ZN(n1000) );
  INV_X1 U1090 ( .A(KEYINPUT55), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(G29), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1035) );
  XNOR2_X1 U1094 ( .A(n1004), .B(G1956), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT119), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1024) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1022) );
  XNOR2_X1 U1099 ( .A(G1348), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(G1971), .A2(G303), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT120), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G1341), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT121), .B(n1025), .ZN(n1031) );
  XNOR2_X1 U1110 ( .A(G1966), .B(G168), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(n1026), .B(KEYINPUT118), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT57), .B(n1029), .Z(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(KEYINPUT56), .B(G16), .Z(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(n1036), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
  INV_X1 U1120 ( .A(G171), .ZN(G301) );
endmodule

