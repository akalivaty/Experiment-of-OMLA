

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795;

  NAND2_X1 U378 ( .A1(n574), .A2(n570), .ZN(n713) );
  XNOR2_X1 U379 ( .A(n629), .B(n374), .ZN(n618) );
  OR2_X2 U380 ( .A1(n688), .A2(G902), .ZN(n484) );
  XNOR2_X2 U381 ( .A(n637), .B(n636), .ZN(n730) );
  NAND2_X1 U382 ( .A1(n357), .A2(n563), .ZN(n586) );
  INV_X1 U383 ( .A(n619), .ZN(n357) );
  INV_X1 U384 ( .A(KEYINPUT35), .ZN(n445) );
  NAND2_X1 U385 ( .A1(n429), .A2(n427), .ZN(n637) );
  AND2_X1 U386 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U387 ( .A1(n432), .A2(n635), .ZN(n431) );
  AND2_X1 U388 ( .A1(n592), .A2(n728), .ZN(n392) );
  NAND2_X1 U389 ( .A1(n405), .A2(n422), .ZN(n687) );
  AND2_X1 U390 ( .A1(n402), .A2(n401), .ZN(n405) );
  NAND2_X1 U391 ( .A1(n378), .A2(n377), .ZN(n383) );
  NOR2_X1 U392 ( .A1(n381), .A2(n379), .ZN(n378) );
  INV_X1 U393 ( .A(n457), .ZN(n399) );
  NAND2_X1 U394 ( .A1(n572), .A2(n610), .ZN(n457) );
  OR2_X1 U395 ( .A1(n722), .A2(n684), .ZN(n580) );
  NOR2_X1 U396 ( .A1(n416), .A2(n415), .ZN(n519) );
  NOR2_X1 U397 ( .A1(n586), .A2(n375), .ZN(n397) );
  INV_X1 U398 ( .A(n744), .ZN(n356) );
  OR2_X1 U399 ( .A1(n437), .A2(n441), .ZN(n590) );
  OR2_X1 U400 ( .A1(n657), .A2(n650), .ZN(n537) );
  XNOR2_X1 U401 ( .A(n785), .B(n476), .ZN(n515) );
  XNOR2_X1 U402 ( .A(n473), .B(n551), .ZN(n527) );
  XNOR2_X1 U403 ( .A(n472), .B(KEYINPUT4), .ZN(n473) );
  XNOR2_X1 U404 ( .A(G119), .B(G116), .ZN(n479) );
  XNOR2_X1 U405 ( .A(n390), .B(n593), .ZN(n598) );
  XNOR2_X1 U406 ( .A(n521), .B(n493), .ZN(n542) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n493) );
  XNOR2_X1 U408 ( .A(n527), .B(n475), .ZN(n785) );
  XNOR2_X1 U409 ( .A(KEYINPUT71), .B(G134), .ZN(n474) );
  BUF_X1 U410 ( .A(n564), .Z(n629) );
  NAND2_X1 U411 ( .A1(n598), .A2(n424), .ZN(n423) );
  NOR2_X1 U412 ( .A1(n679), .A2(n467), .ZN(n424) );
  NAND2_X1 U413 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X1 U414 ( .A(n590), .B(KEYINPUT1), .ZN(n600) );
  XNOR2_X1 U415 ( .A(KEYINPUT5), .B(G137), .ZN(n477) );
  XNOR2_X1 U416 ( .A(n436), .B(n548), .ZN(n667) );
  XNOR2_X1 U417 ( .A(n543), .B(n365), .ZN(n436) );
  NAND2_X1 U418 ( .A1(n577), .A2(n373), .ZN(n376) );
  BUF_X1 U419 ( .A(n600), .Z(n632) );
  NAND2_X1 U420 ( .A1(n399), .A2(n582), .ZN(n406) );
  XNOR2_X1 U421 ( .A(n581), .B(KEYINPUT81), .ZN(n582) );
  NOR2_X1 U422 ( .A1(n585), .A2(KEYINPUT30), .ZN(n420) );
  XNOR2_X1 U423 ( .A(n498), .B(n497), .ZN(n550) );
  XOR2_X1 U424 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n497) );
  XNOR2_X1 U425 ( .A(n496), .B(n495), .ZN(n498) );
  INV_X1 U426 ( .A(KEYINPUT69), .ZN(n495) );
  NAND2_X1 U427 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U428 ( .A(n569), .B(n568), .ZN(n391) );
  NAND2_X1 U429 ( .A1(n453), .A2(n612), .ZN(n382) );
  NAND2_X1 U430 ( .A1(n385), .A2(n446), .ZN(n380) );
  NAND2_X1 U431 ( .A1(n600), .A2(n356), .ZN(n627) );
  XNOR2_X1 U432 ( .A(KEYINPUT16), .B(G122), .ZN(n528) );
  XNOR2_X1 U433 ( .A(G128), .B(G119), .ZN(n499) );
  XNOR2_X1 U434 ( .A(n542), .B(n494), .ZN(n784) );
  XNOR2_X1 U435 ( .A(n464), .B(n463), .ZN(n529) );
  XNOR2_X1 U436 ( .A(G107), .B(G104), .ZN(n464) );
  XNOR2_X1 U437 ( .A(KEYINPUT83), .B(G110), .ZN(n463) );
  XOR2_X1 U438 ( .A(G137), .B(G140), .Z(n511) );
  AND2_X1 U439 ( .A1(n393), .A2(n590), .ZN(n572) );
  AND2_X1 U440 ( .A1(n425), .A2(n395), .ZN(n394) );
  NAND2_X1 U441 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U442 ( .A1(n459), .A2(n358), .ZN(n469) );
  XNOR2_X1 U443 ( .A(n555), .B(G478), .ZN(n573) );
  XNOR2_X1 U444 ( .A(n549), .B(n471), .ZN(n571) );
  XNOR2_X1 U445 ( .A(n444), .B(KEYINPUT32), .ZN(n384) );
  NOR2_X1 U446 ( .A1(n622), .A2(n363), .ZN(n444) );
  NAND2_X1 U447 ( .A1(n632), .A2(n357), .ZN(n400) );
  AND2_X1 U448 ( .A1(n456), .A2(n454), .ZN(n578) );
  XNOR2_X1 U449 ( .A(n455), .B(KEYINPUT91), .ZN(n454) );
  NAND2_X1 U450 ( .A1(n457), .A2(KEYINPUT47), .ZN(n456) );
  NOR2_X1 U451 ( .A1(n580), .A2(n579), .ZN(n455) );
  INV_X1 U452 ( .A(KEYINPUT104), .ZN(n448) );
  NOR2_X1 U453 ( .A1(n631), .A2(n737), .ZN(n449) );
  XNOR2_X1 U454 ( .A(KEYINPUT85), .B(n361), .ZN(n545) );
  INV_X1 U455 ( .A(KEYINPUT76), .ZN(n433) );
  INV_X1 U456 ( .A(n517), .ZN(n440) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  INV_X1 U458 ( .A(G237), .ZN(n485) );
  XNOR2_X1 U459 ( .A(G113), .B(KEYINPUT74), .ZN(n480) );
  XNOR2_X1 U460 ( .A(KEYINPUT70), .B(G131), .ZN(n544) );
  XNOR2_X1 U461 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n541) );
  XNOR2_X1 U462 ( .A(G143), .B(G113), .ZN(n539) );
  XOR2_X1 U463 ( .A(G122), .B(G104), .Z(n540) );
  XNOR2_X1 U464 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n523) );
  XNOR2_X1 U465 ( .A(n627), .B(n601), .ZN(n602) );
  NOR2_X1 U466 ( .A1(n418), .A2(n560), .ZN(n417) );
  XNOR2_X1 U467 ( .A(G134), .B(G116), .ZN(n554) );
  XNOR2_X1 U468 ( .A(n553), .B(n368), .ZN(n409) );
  XOR2_X1 U469 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n553) );
  AND2_X1 U470 ( .A1(n426), .A2(n652), .ZN(n653) );
  INV_X1 U471 ( .A(KEYINPUT40), .ZN(n458) );
  NAND2_X1 U472 ( .A1(n380), .A2(n364), .ZN(n379) );
  NOR2_X1 U473 ( .A1(n765), .A2(n382), .ZN(n381) );
  INV_X1 U474 ( .A(KEYINPUT0), .ZN(n386) );
  NAND2_X1 U475 ( .A1(n452), .A2(n398), .ZN(n752) );
  INV_X1 U476 ( .A(n632), .ZN(n745) );
  XNOR2_X1 U477 ( .A(n689), .B(KEYINPUT62), .ZN(n690) );
  XNOR2_X1 U478 ( .A(n462), .B(n461), .ZN(n695) );
  XNOR2_X1 U479 ( .A(n784), .B(n503), .ZN(n462) );
  XNOR2_X1 U480 ( .A(n410), .B(n407), .ZN(n701) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U482 ( .A(n411), .B(n552), .ZN(n410) );
  XNOR2_X1 U483 ( .A(n554), .B(KEYINPUT7), .ZN(n408) );
  XNOR2_X1 U484 ( .A(n667), .B(n666), .ZN(n668) );
  BUF_X1 U485 ( .A(n700), .Z(n705) );
  XNOR2_X1 U486 ( .A(n515), .B(n514), .ZN(n707) );
  XNOR2_X1 U487 ( .A(n657), .B(n659), .ZN(n660) );
  INV_X2 U488 ( .A(G953), .ZN(n788) );
  NAND2_X1 U489 ( .A1(n413), .A2(n572), .ZN(n567) );
  INV_X1 U490 ( .A(n764), .ZN(n413) );
  NOR2_X1 U491 ( .A1(n599), .A2(n718), .ZN(n679) );
  XNOR2_X1 U492 ( .A(n450), .B(KEYINPUT31), .ZN(n723) );
  NAND2_X1 U493 ( .A1(n453), .A2(n451), .ZN(n450) );
  INV_X1 U494 ( .A(n752), .ZN(n451) );
  XNOR2_X1 U495 ( .A(n412), .B(KEYINPUT103), .ZN(n722) );
  XNOR2_X1 U496 ( .A(n387), .B(KEYINPUT106), .ZN(n680) );
  NAND2_X1 U497 ( .A1(n633), .A2(n389), .ZN(n388) );
  INV_X1 U498 ( .A(n618), .ZN(n389) );
  XNOR2_X1 U499 ( .A(n384), .B(n681), .ZN(G21) );
  NOR2_X1 U500 ( .A1(n556), .A2(n373), .ZN(n358) );
  AND2_X1 U501 ( .A1(n376), .A2(n372), .ZN(n359) );
  AND2_X1 U502 ( .A1(n470), .A2(n684), .ZN(n360) );
  OR2_X1 U503 ( .A1(G953), .A2(G237), .ZN(n361) );
  XOR2_X1 U504 ( .A(n508), .B(n507), .Z(n362) );
  INV_X1 U505 ( .A(n747), .ZN(n414) );
  OR2_X1 U506 ( .A1(n618), .A2(n400), .ZN(n363) );
  XOR2_X1 U507 ( .A(n614), .B(KEYINPUT88), .Z(n364) );
  XOR2_X1 U508 ( .A(n540), .B(n539), .Z(n365) );
  XOR2_X1 U509 ( .A(n482), .B(n530), .Z(n366) );
  AND2_X1 U510 ( .A1(n615), .A2(n414), .ZN(n367) );
  XOR2_X1 U511 ( .A(G107), .B(G122), .Z(n368) );
  AND2_X1 U512 ( .A1(n466), .A2(n587), .ZN(n369) );
  INV_X1 U513 ( .A(G902), .ZN(n439) );
  AND2_X1 U514 ( .A1(n630), .A2(n629), .ZN(n370) );
  AND2_X1 U515 ( .A1(n358), .A2(KEYINPUT40), .ZN(n371) );
  AND2_X1 U516 ( .A1(n360), .A2(n458), .ZN(n372) );
  XNOR2_X1 U517 ( .A(KEYINPUT77), .B(KEYINPUT39), .ZN(n373) );
  XOR2_X1 U518 ( .A(KEYINPUT105), .B(KEYINPUT6), .Z(n374) );
  XNOR2_X1 U519 ( .A(n565), .B(KEYINPUT28), .ZN(n375) );
  NAND2_X1 U520 ( .A1(n376), .A2(n360), .ZN(n403) );
  NAND2_X1 U521 ( .A1(n468), .A2(n376), .ZN(n599) );
  NAND2_X1 U522 ( .A1(n765), .A2(n446), .ZN(n377) );
  XNOR2_X2 U523 ( .A(n605), .B(n604), .ZN(n765) );
  XNOR2_X2 U524 ( .A(n383), .B(n445), .ZN(n686) );
  NAND2_X1 U525 ( .A1(n618), .A2(n369), .ZN(n594) );
  NOR2_X1 U526 ( .A1(n384), .A2(n677), .ZN(n625) );
  AND2_X1 U527 ( .A1(n453), .A2(n370), .ZN(n712) );
  INV_X1 U528 ( .A(n453), .ZN(n385) );
  XNOR2_X2 U529 ( .A(n611), .B(n386), .ZN(n453) );
  OR2_X1 U530 ( .A1(n622), .A2(n388), .ZN(n387) );
  NAND2_X1 U531 ( .A1(n396), .A2(n394), .ZN(n393) );
  NAND2_X1 U532 ( .A1(n586), .A2(n375), .ZN(n395) );
  INV_X1 U533 ( .A(n629), .ZN(n398) );
  NAND2_X1 U534 ( .A1(n399), .A2(n722), .ZN(n673) );
  NAND2_X1 U535 ( .A1(n399), .A2(n684), .ZN(n685) );
  NAND2_X1 U536 ( .A1(n459), .A2(n371), .ZN(n401) );
  NAND2_X1 U537 ( .A1(n403), .A2(KEYINPUT40), .ZN(n402) );
  XNOR2_X2 U538 ( .A(n404), .B(KEYINPUT86), .ZN(n577) );
  NAND2_X1 U539 ( .A1(n518), .A2(n519), .ZN(n404) );
  NAND2_X1 U540 ( .A1(n421), .A2(n420), .ZN(n419) );
  XNOR2_X1 U541 ( .A(n406), .B(KEYINPUT80), .ZN(n583) );
  NAND2_X1 U542 ( .A1(n550), .A2(G217), .ZN(n411) );
  INV_X1 U543 ( .A(n573), .ZN(n570) );
  NAND2_X1 U544 ( .A1(n571), .A2(n573), .ZN(n412) );
  NAND2_X1 U545 ( .A1(n619), .A2(n414), .ZN(n744) );
  XNOR2_X2 U546 ( .A(n460), .B(n362), .ZN(n619) );
  AND2_X1 U547 ( .A1(n564), .A2(KEYINPUT30), .ZN(n415) );
  NAND2_X1 U548 ( .A1(n419), .A2(n417), .ZN(n416) );
  AND2_X1 U549 ( .A1(n585), .A2(KEYINPUT30), .ZN(n418) );
  INV_X1 U550 ( .A(n564), .ZN(n421) );
  XNOR2_X2 U551 ( .A(n484), .B(n483), .ZN(n564) );
  NAND2_X1 U552 ( .A1(n359), .A2(n469), .ZN(n422) );
  NAND2_X1 U553 ( .A1(n687), .A2(n676), .ZN(n569) );
  XNOR2_X2 U554 ( .A(n423), .B(KEYINPUT93), .ZN(n731) );
  NAND2_X1 U555 ( .A1(n564), .A2(n375), .ZN(n425) );
  NAND2_X1 U556 ( .A1(n734), .A2(n426), .ZN(n763) );
  NAND2_X1 U557 ( .A1(n648), .A2(n730), .ZN(n426) );
  XNOR2_X1 U558 ( .A(n623), .B(n433), .ZN(n428) );
  NAND2_X1 U559 ( .A1(n428), .A2(n626), .ZN(n427) );
  XNOR2_X1 U560 ( .A(n434), .B(KEYINPUT107), .ZN(n430) );
  NAND2_X1 U561 ( .A1(n626), .A2(KEYINPUT44), .ZN(n432) );
  NAND2_X1 U562 ( .A1(n447), .A2(n680), .ZN(n434) );
  XNOR2_X1 U563 ( .A(n435), .B(KEYINPUT79), .ZN(n592) );
  NAND2_X1 U564 ( .A1(n583), .A2(n584), .ZN(n435) );
  NAND2_X1 U565 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U566 ( .A(n577), .ZN(n459) );
  NOR2_X1 U567 ( .A1(n707), .A2(n438), .ZN(n437) );
  NAND2_X1 U568 ( .A1(n517), .A2(G902), .ZN(n442) );
  NAND2_X1 U569 ( .A1(n707), .A2(n517), .ZN(n443) );
  NAND2_X1 U570 ( .A1(n686), .A2(n625), .ZN(n623) );
  INV_X1 U571 ( .A(n612), .ZN(n446) );
  XNOR2_X1 U572 ( .A(n449), .B(n448), .ZN(n447) );
  INV_X1 U573 ( .A(n627), .ZN(n452) );
  INV_X1 U574 ( .A(n580), .ZN(n737) );
  NAND2_X1 U575 ( .A1(n695), .A2(n439), .ZN(n460) );
  XNOR2_X1 U576 ( .A(n502), .B(KEYINPUT100), .ZN(n461) );
  INV_X1 U577 ( .A(n575), .ZN(n596) );
  NAND2_X1 U578 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X2 U579 ( .A(n465), .B(KEYINPUT19), .ZN(n610) );
  NAND2_X1 U580 ( .A1(n575), .A2(n466), .ZN(n465) );
  INV_X1 U581 ( .A(n585), .ZN(n466) );
  NAND2_X1 U582 ( .A1(n598), .A2(n678), .ZN(n647) );
  INV_X1 U583 ( .A(n678), .ZN(n467) );
  AND2_X1 U584 ( .A1(n469), .A2(n470), .ZN(n468) );
  NAND2_X1 U585 ( .A1(n556), .A2(n373), .ZN(n470) );
  XNOR2_X1 U586 ( .A(KEYINPUT13), .B(G475), .ZN(n471) );
  INV_X1 U587 ( .A(KEYINPUT46), .ZN(n568) );
  INV_X1 U588 ( .A(KEYINPUT108), .ZN(n601) );
  INV_X1 U589 ( .A(n511), .ZN(n494) );
  XNOR2_X1 U590 ( .A(n486), .B(KEYINPUT99), .ZN(n585) );
  BUF_X1 U591 ( .A(n731), .Z(n787) );
  BUF_X1 U592 ( .A(n730), .Z(n771) );
  INV_X1 U593 ( .A(KEYINPUT60), .ZN(n671) );
  XNOR2_X2 U594 ( .A(G128), .B(KEYINPUT64), .ZN(n472) );
  XNOR2_X1 U595 ( .A(KEYINPUT65), .B(G143), .ZN(n551) );
  XNOR2_X1 U596 ( .A(n544), .B(n474), .ZN(n475) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(G101), .ZN(n520) );
  XNOR2_X1 U598 ( .A(n520), .B(G146), .ZN(n476) );
  NAND2_X1 U599 ( .A1(n545), .A2(G210), .ZN(n478) );
  XNOR2_X1 U600 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U601 ( .A(n479), .B(KEYINPUT3), .ZN(n481) );
  XNOR2_X1 U602 ( .A(n481), .B(n480), .ZN(n530) );
  XNOR2_X1 U603 ( .A(n515), .B(n366), .ZN(n688) );
  INV_X1 U604 ( .A(G472), .ZN(n483) );
  NAND2_X1 U605 ( .A1(n439), .A2(n485), .ZN(n533) );
  NAND2_X1 U606 ( .A1(n533), .A2(G214), .ZN(n486) );
  NAND2_X1 U607 ( .A1(G234), .A2(G237), .ZN(n487) );
  XNOR2_X1 U608 ( .A(n487), .B(KEYINPUT14), .ZN(n735) );
  NOR2_X1 U609 ( .A1(G902), .A2(n788), .ZN(n489) );
  NOR2_X1 U610 ( .A1(G953), .A2(G952), .ZN(n488) );
  NOR2_X1 U611 ( .A1(n489), .A2(n488), .ZN(n490) );
  AND2_X1 U612 ( .A1(n735), .A2(n490), .ZN(n606) );
  NAND2_X1 U613 ( .A1(G953), .A2(G900), .ZN(n491) );
  NAND2_X1 U614 ( .A1(n606), .A2(n491), .ZN(n560) );
  INV_X2 U615 ( .A(G146), .ZN(n492) );
  XNOR2_X2 U616 ( .A(n492), .B(G125), .ZN(n521) );
  NAND2_X1 U617 ( .A1(G234), .A2(n788), .ZN(n496) );
  NAND2_X1 U618 ( .A1(n550), .A2(G221), .ZN(n503) );
  XOR2_X1 U619 ( .A(KEYINPUT23), .B(G110), .Z(n500) );
  XNOR2_X1 U620 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U621 ( .A(n501), .B(KEYINPUT24), .ZN(n502) );
  XOR2_X1 U622 ( .A(KEYINPUT25), .B(KEYINPUT87), .Z(n506) );
  NAND2_X1 U623 ( .A1(n640), .A2(G234), .ZN(n504) );
  XNOR2_X1 U624 ( .A(n504), .B(KEYINPUT20), .ZN(n509) );
  NAND2_X1 U625 ( .A1(G217), .A2(n509), .ZN(n505) );
  XNOR2_X1 U626 ( .A(n506), .B(n505), .ZN(n508) );
  INV_X1 U627 ( .A(KEYINPUT101), .ZN(n507) );
  NAND2_X1 U628 ( .A1(n509), .A2(G221), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n510), .B(KEYINPUT21), .ZN(n747) );
  NAND2_X1 U630 ( .A1(n788), .A2(G227), .ZN(n512) );
  XNOR2_X1 U631 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U632 ( .A(n529), .B(n513), .ZN(n514) );
  INV_X1 U633 ( .A(KEYINPUT73), .ZN(n516) );
  XNOR2_X1 U634 ( .A(n516), .B(G469), .ZN(n517) );
  NAND2_X1 U635 ( .A1(n356), .A2(n590), .ZN(n628) );
  XNOR2_X1 U636 ( .A(n628), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U637 ( .A(n521), .B(n520), .ZN(n525) );
  NAND2_X1 U638 ( .A1(n788), .A2(G224), .ZN(n522) );
  XNOR2_X1 U639 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U640 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U641 ( .A(n527), .B(n526), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U643 ( .A(n531), .B(n530), .ZN(n778) );
  XNOR2_X1 U644 ( .A(n532), .B(n778), .ZN(n657) );
  INV_X1 U645 ( .A(n640), .ZN(n650) );
  NAND2_X1 U646 ( .A1(n533), .A2(G210), .ZN(n535) );
  INV_X1 U647 ( .A(KEYINPUT98), .ZN(n534) );
  XNOR2_X1 U648 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X2 U649 ( .A(n537), .B(n536), .ZN(n575) );
  XNOR2_X1 U650 ( .A(KEYINPUT82), .B(KEYINPUT38), .ZN(n538) );
  XNOR2_X1 U651 ( .A(n575), .B(n538), .ZN(n556) );
  XNOR2_X1 U652 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U653 ( .A(n544), .B(G140), .ZN(n547) );
  NAND2_X1 U654 ( .A1(n545), .A2(G214), .ZN(n546) );
  XNOR2_X1 U655 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U656 ( .A1(n667), .A2(n439), .ZN(n549) );
  INV_X1 U657 ( .A(n571), .ZN(n574) );
  XNOR2_X1 U658 ( .A(n551), .B(G128), .ZN(n552) );
  NAND2_X1 U659 ( .A1(n701), .A2(n439), .ZN(n555) );
  NAND2_X1 U660 ( .A1(n571), .A2(n570), .ZN(n739) );
  NOR2_X1 U661 ( .A1(n739), .A2(n585), .ZN(n557) );
  INV_X1 U662 ( .A(n556), .ZN(n738) );
  NAND2_X1 U663 ( .A1(n557), .A2(n738), .ZN(n559) );
  XNOR2_X1 U664 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n558) );
  XNOR2_X1 U665 ( .A(n559), .B(n558), .ZN(n764) );
  OR2_X1 U666 ( .A1(n747), .A2(n560), .ZN(n562) );
  INV_X1 U667 ( .A(KEYINPUT72), .ZN(n561) );
  XNOR2_X1 U668 ( .A(n562), .B(n561), .ZN(n563) );
  INV_X1 U669 ( .A(KEYINPUT110), .ZN(n565) );
  XNOR2_X1 U670 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n566) );
  XNOR2_X1 U671 ( .A(n567), .B(n566), .ZN(n676) );
  INV_X1 U672 ( .A(n713), .ZN(n684) );
  AND2_X1 U673 ( .A1(n574), .A2(n573), .ZN(n613) );
  NAND2_X1 U674 ( .A1(n613), .A2(n575), .ZN(n576) );
  OR2_X1 U675 ( .A1(n577), .A2(n576), .ZN(n675) );
  AND2_X2 U676 ( .A1(n578), .A2(n675), .ZN(n584) );
  INV_X1 U677 ( .A(KEYINPUT47), .ZN(n579) );
  NAND2_X1 U678 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U679 ( .A1(n713), .A2(n586), .ZN(n587) );
  OR2_X1 U680 ( .A1(n594), .A2(n596), .ZN(n589) );
  INV_X1 U681 ( .A(KEYINPUT36), .ZN(n588) );
  XNOR2_X1 U682 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n591), .A2(n632), .ZN(n728) );
  INV_X1 U684 ( .A(KEYINPUT48), .ZN(n593) );
  OR2_X1 U685 ( .A1(n594), .A2(n632), .ZN(n595) );
  XNOR2_X1 U686 ( .A(n595), .B(KEYINPUT43), .ZN(n597) );
  NAND2_X1 U687 ( .A1(n597), .A2(n596), .ZN(n678) );
  INV_X1 U688 ( .A(n722), .ZN(n718) );
  XNOR2_X1 U689 ( .A(n731), .B(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U690 ( .A1(n602), .A2(n618), .ZN(n605) );
  XNOR2_X1 U691 ( .A(KEYINPUT96), .B(KEYINPUT33), .ZN(n603) );
  XNOR2_X1 U692 ( .A(n603), .B(KEYINPUT75), .ZN(n604) );
  INV_X1 U693 ( .A(n606), .ZN(n608) );
  AND2_X1 U694 ( .A1(G953), .A2(G898), .ZN(n607) );
  NOR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U696 ( .A(KEYINPUT89), .B(KEYINPUT34), .ZN(n612) );
  INV_X1 U697 ( .A(n613), .ZN(n614) );
  INV_X1 U698 ( .A(n739), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n453), .A2(n367), .ZN(n617) );
  XNOR2_X1 U700 ( .A(KEYINPUT78), .B(KEYINPUT22), .ZN(n616) );
  XNOR2_X1 U701 ( .A(n617), .B(n616), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n619), .A2(n398), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n745), .A2(n620), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n677) );
  AND2_X1 U705 ( .A1(KEYINPUT76), .A2(KEYINPUT44), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U707 ( .A(n628), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n723), .A2(n712), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n357), .ZN(n633) );
  INV_X1 U710 ( .A(n686), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n634), .A2(KEYINPUT44), .ZN(n635) );
  XNOR2_X1 U712 ( .A(KEYINPUT94), .B(KEYINPUT45), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n638), .A2(n730), .ZN(n643) );
  NAND2_X1 U714 ( .A1(KEYINPUT2), .A2(KEYINPUT92), .ZN(n641) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n732) );
  NOR2_X1 U716 ( .A1(n732), .A2(KEYINPUT92), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n649) );
  AND2_X1 U718 ( .A1(n641), .A2(n649), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n654) );
  INV_X1 U720 ( .A(n679), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT90), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  INV_X1 U724 ( .A(n649), .ZN(n651) );
  OR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n656) );
  INV_X1 U727 ( .A(KEYINPUT66), .ZN(n655) );
  XNOR2_X2 U728 ( .A(n656), .B(n655), .ZN(n700) );
  NAND2_X1 U729 ( .A1(n700), .A2(G210), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n658) );
  XOR2_X1 U731 ( .A(n658), .B(KEYINPUT55), .Z(n659) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n663) );
  INV_X1 U733 ( .A(G952), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n662), .A2(G953), .ZN(n698) );
  NAND2_X1 U735 ( .A1(n663), .A2(n698), .ZN(n665) );
  INV_X1 U736 ( .A(KEYINPUT56), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(G51) );
  NAND2_X1 U738 ( .A1(n700), .A2(G475), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT97), .B(KEYINPUT59), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n670), .A2(n698), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G60) );
  XNOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .ZN(n674) );
  XOR2_X1 U744 ( .A(n674), .B(n673), .Z(G30) );
  XNOR2_X1 U745 ( .A(n675), .B(G143), .ZN(G45) );
  XNOR2_X1 U746 ( .A(n676), .B(G137), .ZN(G39) );
  XOR2_X1 U747 ( .A(G110), .B(n677), .Z(G12) );
  XNOR2_X1 U748 ( .A(n678), .B(G140), .ZN(G42) );
  XOR2_X1 U749 ( .A(G134), .B(n679), .Z(G36) );
  XNOR2_X1 U750 ( .A(n680), .B(G101), .ZN(G3) );
  XNOR2_X1 U751 ( .A(G119), .B(KEYINPUT127), .ZN(n681) );
  XNOR2_X1 U752 ( .A(G113), .B(KEYINPUT115), .ZN(n683) );
  NAND2_X1 U753 ( .A1(n723), .A2(n684), .ZN(n682) );
  XOR2_X1 U754 ( .A(n683), .B(n682), .Z(G15) );
  XNOR2_X1 U755 ( .A(n685), .B(G146), .ZN(G48) );
  XNOR2_X1 U756 ( .A(n686), .B(G122), .ZN(G24) );
  XNOR2_X1 U757 ( .A(n687), .B(G131), .ZN(G33) );
  NAND2_X1 U758 ( .A1(n700), .A2(G472), .ZN(n691) );
  INV_X1 U759 ( .A(n688), .ZN(n689) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n692), .A2(n698), .ZN(n694) );
  XOR2_X1 U762 ( .A(KEYINPUT95), .B(KEYINPUT63), .Z(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(G57) );
  NAND2_X1 U764 ( .A1(n705), .A2(G217), .ZN(n697) );
  INV_X1 U765 ( .A(n695), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(n699) );
  INV_X1 U767 ( .A(n698), .ZN(n710) );
  NOR2_X1 U768 ( .A1(n699), .A2(n710), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n705), .A2(G478), .ZN(n703) );
  XOR2_X1 U770 ( .A(n701), .B(KEYINPUT122), .Z(n702) );
  XNOR2_X1 U771 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U772 ( .A1(n704), .A2(n710), .ZN(G63) );
  NAND2_X1 U773 ( .A1(n705), .A2(G469), .ZN(n709) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XNOR2_X1 U775 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(G54) );
  INV_X1 U778 ( .A(n712), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n719), .A2(n713), .ZN(n715) );
  XNOR2_X1 U780 ( .A(G104), .B(KEYINPUT113), .ZN(n714) );
  XNOR2_X1 U781 ( .A(n715), .B(n714), .ZN(G6) );
  XOR2_X1 U782 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n717) );
  XNOR2_X1 U783 ( .A(G107), .B(KEYINPUT27), .ZN(n716) );
  XNOR2_X1 U784 ( .A(n717), .B(n716), .ZN(n721) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U786 ( .A(n721), .B(n720), .Z(G9) );
  XNOR2_X1 U787 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n725) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U789 ( .A(n725), .B(n724), .Z(n726) );
  XNOR2_X1 U790 ( .A(G116), .B(n726), .ZN(G18) );
  XOR2_X1 U791 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n727) );
  XNOR2_X1 U792 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U793 ( .A(G125), .B(n729), .ZN(G27) );
  NAND2_X1 U794 ( .A1(n771), .A2(n787), .ZN(n733) );
  NAND2_X1 U795 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U796 ( .A1(G952), .A2(n735), .ZN(n760) );
  NAND2_X1 U797 ( .A1(n738), .A2(n466), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n742) );
  NOR2_X1 U799 ( .A1(n738), .A2(n466), .ZN(n740) );
  NOR2_X1 U800 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n765), .A2(n743), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U804 ( .A(n746), .B(KEYINPUT50), .ZN(n751) );
  NAND2_X1 U805 ( .A1(n357), .A2(n747), .ZN(n748) );
  XNOR2_X1 U806 ( .A(n748), .B(KEYINPUT49), .ZN(n749) );
  NOR2_X1 U807 ( .A1(n749), .A2(n398), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U809 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U810 ( .A(n754), .B(KEYINPUT51), .ZN(n755) );
  NOR2_X1 U811 ( .A1(n755), .A2(n764), .ZN(n756) );
  OR2_X1 U812 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U813 ( .A(KEYINPUT52), .B(n758), .Z(n759) );
  NOR2_X1 U814 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U815 ( .A(n761), .B(KEYINPUT119), .ZN(n762) );
  NAND2_X1 U816 ( .A1(n763), .A2(n762), .ZN(n768) );
  NOR2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n766), .B(KEYINPUT120), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U820 ( .A1(n788), .A2(n769), .ZN(n770) );
  XOR2_X1 U821 ( .A(KEYINPUT53), .B(n770), .Z(G75) );
  INV_X1 U822 ( .A(n771), .ZN(n772) );
  NOR2_X1 U823 ( .A1(n772), .A2(G953), .ZN(n777) );
  NAND2_X1 U824 ( .A1(G953), .A2(G224), .ZN(n773) );
  XNOR2_X1 U825 ( .A(KEYINPUT61), .B(n773), .ZN(n774) );
  NAND2_X1 U826 ( .A1(n774), .A2(G898), .ZN(n775) );
  XNOR2_X1 U827 ( .A(n775), .B(KEYINPUT123), .ZN(n776) );
  NOR2_X1 U828 ( .A1(n777), .A2(n776), .ZN(n783) );
  XOR2_X1 U829 ( .A(G101), .B(n778), .Z(n780) );
  NOR2_X1 U830 ( .A1(G898), .A2(n788), .ZN(n779) );
  NOR2_X1 U831 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U832 ( .A(KEYINPUT124), .B(n781), .Z(n782) );
  XNOR2_X1 U833 ( .A(n783), .B(n782), .ZN(G69) );
  XNOR2_X1 U834 ( .A(n784), .B(KEYINPUT125), .ZN(n786) );
  XNOR2_X1 U835 ( .A(n785), .B(n786), .ZN(n791) );
  XOR2_X1 U836 ( .A(n791), .B(n787), .Z(n789) );
  NAND2_X1 U837 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U838 ( .A(n790), .B(KEYINPUT126), .ZN(n795) );
  XNOR2_X1 U839 ( .A(G227), .B(n791), .ZN(n792) );
  NAND2_X1 U840 ( .A1(n792), .A2(G900), .ZN(n793) );
  NAND2_X1 U841 ( .A1(n793), .A2(G953), .ZN(n794) );
  NAND2_X1 U842 ( .A1(n795), .A2(n794), .ZN(G72) );
endmodule

