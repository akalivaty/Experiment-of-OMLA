//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT84), .Z(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n207), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(G155gat), .B2(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT81), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n206), .A2(new_n207), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(KEYINPUT80), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n216), .ZN(new_n226));
  INV_X1    g025(.A(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G211gat), .B(G218gat), .Z(new_n232));
  INV_X1    g031(.A(G197gat), .ZN(new_n233));
  INV_X1    g032(.A(G204gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT22), .ZN(new_n237));
  NAND2_X1  g036(.A1(G211gat), .A2(G218gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n235), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n232), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n237), .ZN(new_n242));
  INV_X1    g041(.A(new_n236), .ZN(new_n243));
  NOR2_X1   g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT73), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n247), .A3(KEYINPUT74), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(KEYINPUT75), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n241), .A2(new_n247), .A3(KEYINPUT74), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT74), .B1(new_n241), .B2(new_n247), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT86), .B1(new_n248), .B2(KEYINPUT29), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT86), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n241), .A2(new_n247), .A3(new_n259), .A4(new_n230), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n222), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n221), .A2(new_n228), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n257), .A2(new_n263), .A3(G228gat), .A4(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G228gat), .A2(G233gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n215), .A2(new_n220), .B1(new_n226), .B2(new_n227), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n239), .A2(new_n232), .A3(KEYINPUT85), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n245), .B1(new_n268), .B2(new_n246), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n267), .A2(new_n269), .B1(new_n268), .B2(new_n246), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n230), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n271), .B2(new_n222), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n229), .A2(new_n230), .B1(new_n251), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n265), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G22gat), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n264), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n203), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n264), .A2(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G22gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n203), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT31), .B(G50gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n278), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n278), .B2(new_n283), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G85gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT87), .Z(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(G113gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G120gat), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n294), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n298), .B1(new_n297), .B2(new_n304), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT4), .B1(new_n308), .B2(new_n262), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n305), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n266), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(KEYINPUT82), .A3(new_n305), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n306), .B2(new_n307), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .A4(new_n229), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n293), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT39), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n292), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n320), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT39), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n318), .A2(new_n316), .A3(new_n262), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n311), .A2(new_n266), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n293), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT40), .B(new_n322), .C1(new_n324), .C2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n319), .A3(KEYINPUT5), .A4(new_n293), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n314), .A2(new_n293), .A3(new_n319), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(new_n293), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n331), .B(new_n292), .C1(new_n332), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n327), .B(KEYINPUT88), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT39), .A3(new_n323), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT40), .B1(new_n340), .B2(new_n322), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT27), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT27), .B(G183gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n345), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n344), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n346), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT28), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT66), .B(G183gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n360), .B2(KEYINPUT27), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT67), .B(new_n359), .C1(new_n361), .C2(new_n347), .ZN(new_n362));
  INV_X1    g161(.A(G169gat), .ZN(new_n363));
  INV_X1    g162(.A(G176gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT68), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n365), .A2(KEYINPUT26), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n365), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n366), .A2(new_n367), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n356), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT23), .B1(new_n363), .B2(new_n364), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n364), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G183gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(KEYINPUT24), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n378), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n372), .B(new_n376), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n373), .B2(new_n364), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n360), .A2(G190gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n372), .B(new_n386), .C1(new_n387), .C2(new_n380), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT29), .B1(new_n369), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT78), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n369), .A2(new_n389), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n391), .B(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n254), .A2(new_n255), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n256), .A2(new_n252), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n396), .B1(new_n395), .B2(new_n230), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n391), .B1(new_n369), .B2(new_n389), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n395), .A2(new_n392), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n390), .B2(new_n396), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n407), .B2(new_n401), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G8gat), .B(G36gat), .Z(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n399), .B(new_n412), .C1(new_n405), .C2(new_n408), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n343), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n343), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n342), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT38), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n409), .B2(KEYINPUT37), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n421), .A2(KEYINPUT90), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(new_n412), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n331), .B1(new_n332), .B2(new_n336), .ZN(new_n431));
  INV_X1    g230(.A(new_n291), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n291), .B(new_n331), .C1(new_n332), .C2(new_n336), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n433), .A2(new_n337), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n437));
  INV_X1    g236(.A(new_n398), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT89), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n407), .A2(new_n401), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(KEYINPUT89), .A3(new_n438), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n420), .B(new_n413), .C1(new_n409), .C2(KEYINPUT37), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n436), .B(new_n415), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n287), .B(new_n419), .C1(new_n428), .C2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(G15gat), .B(G43gat), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT71), .ZN(new_n448));
  XOR2_X1   g247(.A(G71gat), .B(G99gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n395), .A2(new_n311), .ZN(new_n451));
  INV_X1    g250(.A(G227gat), .ZN(new_n452));
  INV_X1    g251(.A(G233gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n308), .A2(new_n369), .A3(new_n389), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(KEYINPUT32), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n456), .B(KEYINPUT32), .C1(new_n458), .C2(new_n450), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n451), .A2(new_n455), .ZN(new_n464));
  INV_X1    g263(.A(new_n454), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n463), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n463), .B2(KEYINPUT72), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT36), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n470), .A2(new_n461), .A3(new_n462), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n461), .B2(new_n462), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n285), .A2(new_n286), .ZN(new_n479));
  INV_X1    g278(.A(new_n416), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n433), .A2(new_n434), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n435), .A2(new_n430), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n483), .A3(new_n417), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n478), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n446), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n472), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n463), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n487), .B(new_n488), .C1(new_n285), .C2(new_n286), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT35), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n416), .A2(new_n418), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n475), .A2(new_n476), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n287), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n275), .A2(G15gat), .ZN(new_n497));
  INV_X1    g296(.A(G15gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G22gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT94), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT95), .B1(new_n501), .B2(new_n504), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n502), .A2(new_n503), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n509), .A2(G8gat), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n513), .A2(new_n514), .B1(new_n506), .B2(new_n505), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(G1gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G57gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G64gat), .ZN(new_n529));
  INV_X1    g328(.A(G64gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G57gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G71gat), .B(G78gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n526), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT21), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT102), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n536), .A2(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n545), .B(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT101), .B(KEYINPUT19), .Z(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n556), .A3(new_n550), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT14), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(KEYINPUT92), .A2(G29gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(KEYINPUT92), .A2(G29gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(G43gat), .ZN(new_n573));
  INV_X1    g372(.A(G50gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G43gat), .A2(G50gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT15), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n568), .A2(new_n572), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n563), .B1(new_n569), .B2(new_n570), .ZN(new_n583));
  OAI211_X1 g382(.A(KEYINPUT15), .B(new_n577), .C1(new_n583), .C2(new_n567), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n583), .A2(new_n567), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(KEYINPUT93), .A3(new_n578), .A4(new_n580), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(KEYINPUT105), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT105), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(G85gat), .A3(G92gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT104), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G99gat), .ZN(new_n600));
  INV_X1    g399(.A(G106gat), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT8), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(KEYINPUT104), .ZN(new_n603));
  OR2_X1    g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  NOR3_X1   g405(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n596), .A2(new_n598), .ZN(new_n609));
  AND2_X1   g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT7), .B1(new_n610), .B2(new_n595), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n589), .B(new_n591), .C1(new_n607), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT103), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n588), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n614), .A2(new_n607), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n618), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT106), .ZN(new_n629));
  INV_X1    g428(.A(new_n624), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n622), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n625), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n628), .B(KEYINPUT106), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n625), .B2(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n527), .A2(new_n535), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n614), .B2(new_n607), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n612), .A2(new_n608), .A3(new_n613), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n606), .B1(new_n599), .B2(new_n605), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n536), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT107), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n638), .A2(new_n645), .A3(new_n642), .A4(new_n639), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n536), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n642), .ZN(new_n655));
  INV_X1    g454(.A(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n650), .B(KEYINPUT108), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n654), .B1(new_n662), .B2(new_n657), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT109), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(KEYINPUT109), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n659), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n561), .A2(new_n636), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n620), .B1(new_n516), .B2(new_n520), .ZN(new_n669));
  OAI21_X1  g468(.A(G8gat), .B1(new_n509), .B2(new_n515), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n518), .A2(new_n517), .A3(new_n519), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n589), .A2(new_n670), .A3(new_n671), .A4(new_n591), .ZN(new_n672));
  NAND2_X1  g471(.A1(G229gat), .A2(G233gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT18), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n669), .A2(new_n672), .A3(KEYINPUT96), .A4(new_n673), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n676), .A2(KEYINPUT97), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n673), .B(KEYINPUT13), .Z(new_n680));
  NOR3_X1   g479(.A1(new_n516), .A2(new_n620), .A3(new_n520), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n588), .B1(new_n670), .B2(new_n671), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n669), .A2(new_n672), .A3(KEYINPUT18), .A4(new_n673), .ZN(new_n684));
  XNOR2_X1  g483(.A(G113gat), .B(G141gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n233), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT11), .B(G169gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT12), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n683), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n679), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT18), .B1(new_n674), .B2(new_n675), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT97), .B1(new_n692), .B2(new_n678), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n683), .A2(new_n684), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n692), .B2(new_n678), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n689), .B(KEYINPUT91), .Z(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI22_X1  g496(.A1(new_n691), .A2(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n692), .A2(new_n678), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT97), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n679), .A3(new_n690), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n692), .A2(new_n678), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n696), .B1(new_n705), .B2(new_n694), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT98), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n668), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n496), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n483), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n514), .ZN(G1324gat));
  INV_X1    g511(.A(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(new_n492), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n517), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT16), .B(G8gat), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n710), .A2(new_n492), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(KEYINPUT42), .B2(new_n717), .ZN(G1325gat));
  NAND2_X1  g518(.A1(new_n478), .A2(KEYINPUT110), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n473), .A2(new_n721), .A3(new_n477), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G15gat), .B1(new_n710), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n493), .A2(new_n498), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n710), .B2(new_n725), .ZN(G1326gat));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n287), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  AOI21_X1  g528(.A(new_n636), .B1(new_n486), .B2(new_n495), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n698), .A2(new_n699), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n704), .A2(new_n706), .A3(KEYINPUT98), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n560), .A3(new_n667), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(new_n483), .A3(new_n571), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT45), .Z(new_n738));
  INV_X1    g537(.A(new_n446), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n484), .A2(new_n479), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n720), .A3(new_n722), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n495), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT44), .B1(new_n742), .B2(new_n635), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(KEYINPUT44), .B2(new_n730), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n560), .A2(new_n667), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n704), .B2(new_n706), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n571), .B1(new_n747), .B2(new_n483), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n738), .A2(new_n748), .ZN(G1328gat));
  OAI21_X1  g548(.A(G36gat), .B1(new_n747), .B2(new_n492), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n736), .A2(G36gat), .A3(new_n492), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1329gat));
  OAI21_X1  g552(.A(G43gat), .B1(new_n747), .B2(new_n723), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n730), .A2(new_n573), .A3(new_n493), .A4(new_n735), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT47), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n755), .C1(new_n757), .C2(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n635), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n287), .A2(new_n574), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n746), .A4(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n730), .B2(new_n735), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n446), .A2(new_n485), .B1(new_n490), .B2(new_n494), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n771), .A2(KEYINPUT113), .A3(new_n636), .A4(new_n734), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n770), .A2(new_n772), .A3(new_n287), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n762), .B(new_n768), .C1(new_n773), .C2(G50gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n765), .A2(new_n766), .A3(new_n746), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n736), .A2(KEYINPUT113), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n730), .A2(new_n769), .A3(new_n735), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n479), .A3(new_n781), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n779), .A2(new_n767), .B1(new_n782), .B2(new_n574), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n776), .B1(new_n783), .B2(KEYINPUT114), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n778), .B2(new_n784), .ZN(G1331gat));
  NOR4_X1   g584(.A1(new_n560), .A2(new_n667), .A3(new_n698), .A4(new_n635), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n742), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n483), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G57gat), .ZN(G1332gat));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n714), .B1(new_n791), .B2(new_n530), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT115), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n530), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1333gat));
  INV_X1    g595(.A(new_n723), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n493), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(G71gat), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n798), .A2(G71gat), .B1(new_n787), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n479), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  INV_X1    g603(.A(new_n763), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n561), .A2(new_n698), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  INV_X1    g607(.A(new_n806), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n763), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g610(.A1(new_n811), .A2(G85gat), .A3(new_n483), .A4(new_n667), .ZN(new_n812));
  INV_X1    g611(.A(G85gat), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n809), .A2(new_n667), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n744), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n788), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n812), .A2(new_n816), .ZN(G1336gat));
  NAND4_X1  g616(.A1(new_n765), .A2(new_n714), .A3(new_n766), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n492), .A2(new_n667), .A3(G92gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n819), .B2(KEYINPUT116), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n822), .B(new_n824), .ZN(G1337gat));
  NOR4_X1   g624(.A1(new_n811), .A2(G99gat), .A3(new_n799), .A4(new_n667), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n600), .B1(new_n815), .B2(new_n797), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(G1338gat));
  NAND4_X1  g627(.A1(new_n765), .A2(new_n479), .A3(new_n766), .A4(new_n814), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n829), .A2(G106gat), .B1(KEYINPUT117), .B2(KEYINPUT53), .ZN(new_n830));
  INV_X1    g629(.A(new_n666), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n658), .B1(new_n831), .B2(new_n664), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n287), .A2(G106gat), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(new_n833), .C1(new_n807), .C2(new_n810), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(G1339gat));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n649), .A2(new_n838), .A3(new_n661), .ZN(new_n839));
  INV_X1    g638(.A(new_n654), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n648), .A2(new_n660), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n647), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n656), .B1(new_n647), .B2(new_n648), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n838), .B1(new_n647), .B2(new_n842), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n651), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n841), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT119), .B1(new_n850), .B2(new_n659), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n660), .B1(new_n647), .B2(new_n648), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n852), .B(new_n654), .C1(new_n853), .C2(new_n838), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n845), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n847), .B1(new_n651), .B2(new_n848), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n658), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n840), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n855), .B2(new_n856), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n852), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n851), .A2(new_n859), .A3(new_n698), .A4(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n681), .A2(new_n682), .A3(new_n680), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n688), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n832), .A2(new_n704), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n635), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n635), .B(new_n867), .C1(new_n691), .C2(new_n693), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n851), .A3(new_n859), .A4(new_n863), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n560), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n668), .A2(new_n698), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n483), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n489), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n492), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n698), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n874), .A2(new_n875), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n287), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT120), .B(new_n479), .C1(new_n874), .C2(new_n875), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n492), .A2(new_n788), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n799), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n708), .A2(new_n300), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n880), .B1(new_n887), .B2(new_n888), .ZN(G1340gat));
  AOI21_X1  g688(.A(G120gat), .B1(new_n879), .B2(new_n832), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n667), .A2(new_n302), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n887), .B2(new_n891), .ZN(G1341gat));
  XNOR2_X1  g691(.A(KEYINPUT69), .B(G127gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n560), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n561), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n887), .A2(new_n894), .B1(new_n895), .B2(new_n893), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n294), .A3(new_n635), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n294), .B1(new_n887), .B2(new_n635), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n797), .A2(new_n886), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n287), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n860), .B1(new_n846), .B2(new_n849), .ZN(new_n904));
  XOR2_X1   g703(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n905));
  OAI211_X1 g704(.A(new_n857), .B(new_n658), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n731), .B2(new_n732), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n832), .A2(new_n704), .A3(new_n867), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n636), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n561), .B1(new_n909), .B2(new_n872), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n668), .A2(new_n698), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n287), .B1(new_n874), .B2(new_n875), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(KEYINPUT57), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n868), .B1(new_n708), .B2(new_n906), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n873), .B1(new_n916), .B2(new_n636), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n875), .B1(new_n917), .B2(new_n561), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT122), .B1(new_n918), .B2(new_n903), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n901), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G141gat), .B1(new_n920), .B2(new_n708), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n723), .A2(new_n479), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n714), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n876), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n733), .A2(new_n204), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  AOI21_X1  g727(.A(KEYINPUT58), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n698), .B(new_n901), .C1(new_n915), .C2(new_n919), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n931), .A2(G141gat), .B1(new_n926), .B2(new_n928), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1344gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n205), .A3(new_n832), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n667), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(KEYINPUT59), .A3(new_n205), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n882), .A2(new_n479), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT57), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n668), .A2(new_n733), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n902), .B(new_n479), .C1(new_n910), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n901), .A2(new_n832), .ZN(new_n943));
  OAI21_X1  g742(.A(G148gat), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n935), .B1(new_n937), .B2(new_n945), .ZN(G1345gat));
  OAI21_X1  g745(.A(G155gat), .B1(new_n920), .B2(new_n560), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n926), .A2(new_n208), .A3(new_n561), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1346gat));
  OAI211_X1 g748(.A(new_n635), .B(new_n901), .C1(new_n915), .C2(new_n919), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G162gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n209), .A3(new_n635), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1347gat));
  AOI21_X1  g756(.A(new_n788), .B1(new_n874), .B2(new_n875), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(new_n714), .A3(new_n877), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n698), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n492), .A2(new_n788), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n493), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n883), .B2(new_n884), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n708), .A2(new_n363), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n959), .B2(new_n832), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n667), .B1(new_n374), .B2(new_n375), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n965), .B2(new_n969), .ZN(G1349gat));
  OAI21_X1  g769(.A(new_n360), .B1(new_n964), .B2(new_n560), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n959), .A2(new_n354), .A3(new_n561), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n346), .A3(new_n635), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n635), .B(new_n963), .C1(new_n883), .C2(new_n884), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n977), .A3(G190gat), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n977), .B1(new_n976), .B2(G190gat), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT61), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n976), .A2(G190gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n984), .B2(new_n978), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n975), .B1(new_n981), .B2(new_n985), .ZN(G1351gat));
  AND2_X1   g785(.A1(new_n939), .A2(new_n941), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n723), .A2(new_n961), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(new_n233), .A3(new_n708), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n922), .A2(new_n492), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n958), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(G197gat), .B1(new_n992), .B2(new_n698), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n990), .A2(new_n993), .ZN(G1352gat));
  NAND3_X1  g793(.A1(new_n992), .A2(new_n234), .A3(new_n832), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT62), .Z(new_n996));
  OAI21_X1  g795(.A(KEYINPUT127), .B1(new_n989), .B2(new_n667), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G204gat), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n667), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(G1353gat));
  INV_X1    g799(.A(new_n992), .ZN(new_n1001));
  OR3_X1    g800(.A1(new_n1001), .A2(G211gat), .A3(new_n560), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n561), .A3(new_n988), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(G218gat), .B1(new_n989), .B2(new_n636), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n636), .A2(G218gat), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n1001), .B2(new_n1009), .ZN(G1355gat));
endmodule


