//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT66), .B(G244), .Z(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G77), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(G50), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n227), .A2(new_n207), .A3(new_n228), .ZN(new_n229));
  NOR4_X1   g0029(.A1(new_n213), .A2(new_n225), .A3(new_n226), .A4(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G303), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n250), .A2(new_n252), .A3(G264), .A4(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n250), .A2(new_n252), .A3(G257), .A4(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT89), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n254), .A2(KEYINPUT89), .A3(new_n255), .A4(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n248), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT5), .B(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n228), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n247), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G270), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n248), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n262), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT90), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT84), .B(G116), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n228), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G283), .ZN(new_n282));
  INV_X1    g0082(.A(G97), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n207), .C1(G33), .C2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n279), .A2(KEYINPUT20), .A3(new_n281), .A4(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n281), .B(new_n284), .C1(new_n277), .C2(new_n207), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n207), .A3(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n249), .A2(G1), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n291), .A2(new_n281), .A3(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(G116), .B1(new_n291), .B2(new_n278), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n275), .A2(new_n276), .A3(G179), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n289), .B2(new_n294), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(KEYINPUT21), .C1(new_n262), .C2(new_n274), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n262), .A2(new_n301), .A3(new_n274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n276), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT91), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n275), .A2(G179), .A3(new_n295), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT90), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT91), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n299), .A4(new_n296), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n295), .A2(G169), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n275), .ZN(new_n312));
  INV_X1    g0112(.A(new_n275), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n295), .B1(new_n313), .B2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n313), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n304), .A2(new_n308), .A3(new_n312), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n266), .A2(G264), .A3(new_n248), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT95), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT3), .B(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G257), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT94), .B(G294), .Z(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n256), .B1(new_n323), .B2(new_n249), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(G250), .A3(new_n256), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT93), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT93), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n320), .B(new_n271), .C1(new_n248), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n271), .A2(new_n318), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n325), .B(KEYINPUT93), .ZN(new_n333));
  INV_X1    g0133(.A(new_n324), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n315), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n293), .A2(G107), .ZN(new_n340));
  INV_X1    g0140(.A(G107), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT25), .B1(new_n291), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n321), .A2(new_n207), .A3(G87), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT22), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n277), .A2(G33), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT23), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n207), .B2(G107), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n341), .A2(KEYINPUT23), .A3(G20), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n349), .A2(new_n207), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT24), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n347), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n345), .B1(new_n358), .B2(new_n281), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n357), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n347), .B2(new_n353), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n281), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n345), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n329), .A2(new_n301), .B1(new_n337), .B2(new_n297), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n317), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n321), .A2(G244), .A3(new_n256), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT83), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n321), .A2(G244), .A3(new_n256), .A4(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n321), .A2(G250), .A3(G1698), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n373), .A2(new_n375), .A3(new_n282), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n336), .ZN(new_n378));
  INV_X1    g0178(.A(G257), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n271), .B1(new_n379), .B2(new_n273), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G20), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT82), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT6), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n386), .A2(new_n283), .A3(G107), .ZN(new_n387));
  XNOR2_X1  g0187(.A(G97), .B(G107), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n385), .B1(new_n207), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n321), .B2(G20), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n251), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT7), .B(new_n207), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n341), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n281), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n291), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(G97), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n293), .B2(G97), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n382), .A2(new_n297), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n380), .B1(new_n336), .B2(new_n377), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n301), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n382), .A2(G200), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(G190), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n397), .A4(new_n400), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT87), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n321), .A2(G244), .A3(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n321), .A2(new_n256), .ZN(new_n411));
  INV_X1    g0211(.A(G238), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n348), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n336), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n270), .A2(new_n265), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n248), .B(G250), .C1(G1), .C2(new_n264), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n301), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n413), .B2(new_n336), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(G169), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g0221(.A(KEYINPUT15), .B(G87), .Z(new_n422));
  INV_X1    g0222(.A(KEYINPUT85), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT15), .B(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT85), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n293), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n398), .A2(new_n422), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n321), .A2(new_n207), .A3(G68), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT19), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n207), .A2(G33), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n283), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G97), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(G33), .A3(G97), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n207), .B1(new_n440), .B2(new_n432), .ZN(new_n441));
  INV_X1    g0241(.A(G87), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(new_n283), .A3(new_n341), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n435), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n281), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n428), .B(new_n430), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n431), .A2(new_n434), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n443), .B1(new_n449), .B2(G20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n429), .B1(new_n451), .B2(new_n281), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT86), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n428), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n421), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n414), .A2(new_n418), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n293), .A2(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n420), .A2(G190), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n457), .A2(new_n452), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n409), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n297), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n453), .B1(new_n452), .B2(new_n428), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n445), .B1(new_n448), .B2(new_n450), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n293), .A2(new_n424), .A3(new_n426), .ZN(new_n466));
  NOR4_X1   g0266(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT86), .A4(new_n429), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n419), .B(new_n463), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT87), .A3(new_n460), .ZN(new_n469));
  AOI211_X1 g0269(.A(KEYINPUT88), .B(new_n408), .C1(new_n462), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT88), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n397), .A2(new_n400), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(G200), .B2(new_n382), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(new_n406), .B1(new_n401), .B2(new_n403), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n471), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n369), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n321), .A2(new_n391), .A3(G20), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT7), .B1(new_n253), .B2(new_n207), .ZN(new_n479));
  OAI21_X1  g0279(.A(G68), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(G58), .A2(G68), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G58), .A2(G68), .ZN(new_n482));
  OAI21_X1  g0282(.A(G20), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT77), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT77), .B(G20), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n383), .A2(G159), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT16), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n445), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n480), .A2(KEYINPUT76), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n202), .B1(new_n392), .B2(new_n395), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT76), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n492), .A2(KEYINPUT16), .A3(new_n495), .A4(new_n488), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT8), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G58), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT69), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n498), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n398), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n504), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT8), .B(G58), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n280), .B(new_n228), .C1(G1), .C2(new_n207), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n505), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n497), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n248), .A3(G274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n248), .A2(new_n517), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n232), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n250), .A2(new_n252), .A3(G226), .A4(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n250), .A2(new_n252), .A3(G223), .A4(new_n256), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n336), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G179), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n516), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(new_n336), .ZN(new_n533));
  INV_X1    g0333(.A(new_n520), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G232), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(new_n315), .A3(new_n519), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n526), .B2(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n392), .A2(new_n395), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n494), .B1(new_n538), .B2(G68), .ZN(new_n539));
  AOI211_X1 g0339(.A(KEYINPUT76), .B(new_n202), .C1(new_n392), .C2(new_n395), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT16), .A4(new_n487), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n490), .B1(new_n493), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n281), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n515), .B(new_n537), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n497), .A2(KEYINPUT79), .A3(new_n515), .A4(new_n537), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(KEYINPUT17), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT80), .A4(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n546), .B2(KEYINPUT17), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n491), .A2(new_n496), .B1(new_n512), .B2(new_n514), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT17), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(KEYINPUT81), .A3(new_n558), .A4(new_n537), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n532), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n519), .B1(new_n520), .B2(new_n412), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n321), .A2(G232), .A3(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G226), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n440), .C1(new_n411), .C2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n567), .B2(new_n336), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT13), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n568), .A2(new_n569), .ZN(new_n572));
  OAI21_X1  g0372(.A(G169), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT14), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(KEYINPUT73), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT73), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n568), .B2(new_n569), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n575), .A2(G179), .A3(new_n577), .A4(new_n570), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n568), .B(new_n569), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(G169), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n290), .A2(G1), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n207), .A2(G68), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT12), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(KEYINPUT75), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n587));
  XOR2_X1   g0387(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g0388(.A(new_n509), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(G68), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G77), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n433), .A2(new_n591), .B1(new_n207), .B2(G68), .ZN(new_n592));
  INV_X1    g0392(.A(G50), .ZN(new_n593));
  INV_X1    g0393(.A(new_n383), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n592), .A2(KEYINPUT74), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n592), .A2(KEYINPUT74), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n281), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT11), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n590), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n582), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n579), .B2(G200), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n575), .A2(G190), .A3(new_n577), .A4(new_n570), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n321), .A2(G222), .A3(new_n256), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n321), .A2(G1698), .ZN(new_n610));
  INV_X1    g0410(.A(G223), .ZN(new_n611));
  OAI221_X1 g0411(.A(new_n609), .B1(new_n215), .B2(new_n321), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n336), .ZN(new_n613));
  INV_X1    g0413(.A(new_n519), .ZN(new_n614));
  XNOR2_X1  g0414(.A(KEYINPUT68), .B(G226), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n534), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT71), .B1(new_n618), .B2(G190), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n330), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g0420(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n621));
  INV_X1    g0421(.A(G150), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n594), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n502), .A2(new_n504), .ZN(new_n624));
  INV_X1    g0424(.A(new_n433), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n445), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n291), .A2(new_n593), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n593), .B2(new_n509), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT9), .ZN(new_n631));
  OR3_X1    g0431(.A1(new_n620), .A2(new_n631), .A3(KEYINPUT10), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT10), .B1(new_n631), .B2(new_n620), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n617), .B2(new_n297), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT70), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n617), .A2(new_n636), .A3(G179), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT70), .B1(new_n618), .B2(new_n301), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n519), .B1(new_n520), .B2(new_n214), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n610), .A2(new_n412), .B1(new_n341), .B2(new_n321), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n253), .A2(new_n232), .A3(G1698), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n336), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(G169), .ZN(new_n645));
  INV_X1    g0445(.A(new_n215), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n646), .A2(new_n398), .B1(new_n509), .B2(new_n591), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(G20), .B1(new_n422), .B2(new_n625), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n594), .B2(new_n507), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n281), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(new_n301), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(G190), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n650), .C1(new_n330), .C2(new_n644), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n608), .A2(new_n634), .A3(new_n639), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n477), .A2(new_n563), .A3(new_n657), .ZN(G372));
  INV_X1    g0458(.A(new_n532), .ZN(new_n659));
  INV_X1    g0459(.A(new_n653), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n603), .B1(new_n606), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n560), .B1(new_n552), .B2(new_n553), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n634), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n639), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n657), .A2(new_n563), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n455), .A2(new_n461), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n475), .A2(new_n667), .A3(new_n360), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n300), .A2(new_n303), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n312), .A3(new_n367), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n455), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  AOI211_X1 g0472(.A(new_n672), .B(new_n404), .C1(new_n462), .C2(new_n469), .ZN(new_n673));
  INV_X1    g0473(.A(new_n404), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT26), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n665), .A2(new_n677), .ZN(G369));
  NAND4_X1  g0478(.A1(new_n306), .A2(new_n299), .A3(new_n296), .A4(new_n312), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n583), .A2(new_n207), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n295), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n317), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT96), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n689), .A2(KEYINPUT96), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n368), .ZN(new_n695));
  INV_X1    g0495(.A(new_n685), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n359), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n367), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n304), .A2(new_n312), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n685), .B1(new_n700), .B2(new_n308), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n365), .A2(new_n366), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n696), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT97), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n707), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n699), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n210), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n206), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n443), .A2(G116), .ZN(new_n714));
  INV_X1    g0514(.A(new_n227), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n713), .A2(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT28), .Z(new_n717));
  NAND2_X1  g0517(.A1(new_n667), .A2(new_n674), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n455), .B1(new_n718), .B2(KEYINPUT26), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n404), .B1(new_n462), .B2(new_n469), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n721), .B2(KEYINPUT26), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n304), .A2(new_n308), .A3(new_n312), .A4(new_n367), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(new_n668), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n696), .C1(new_n722), .C2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n676), .A2(new_n696), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(KEYINPUT29), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n369), .B(new_n696), .C1(new_n470), .C2(new_n476), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n335), .A2(new_n336), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n402), .A2(new_n729), .A3(new_n420), .A4(new_n320), .ZN(new_n730));
  INV_X1    g0530(.A(new_n302), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n402), .A2(G179), .A3(new_n420), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n313), .A3(new_n329), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n732), .B1(new_n730), .B2(new_n731), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n737), .B2(new_n685), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n727), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n717), .B1(new_n743), .B2(G1), .ZN(G364));
  OR2_X1    g0544(.A1(new_n688), .A2(G330), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT98), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n290), .A2(G20), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT99), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n713), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n693), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n750), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n210), .A2(new_n321), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n210), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n711), .A2(new_n321), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n264), .B2(new_n715), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n242), .A2(new_n264), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n228), .B1(G20), .B2(new_n297), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n752), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(new_n301), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n315), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n201), .B1(new_n215), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n207), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n330), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n341), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n774), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(new_n772), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n786));
  XNOR2_X1  g0586(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT103), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n768), .A2(new_n788), .A3(new_n778), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n768), .B2(new_n778), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n787), .B1(G68), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n315), .A2(new_n330), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n779), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n442), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT102), .B1(new_n796), .B2(new_n253), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n796), .A2(KEYINPUT102), .A3(new_n253), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT100), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n768), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n768), .B2(new_n794), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n798), .B1(G50), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n782), .A2(new_n793), .A3(new_n797), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n773), .A2(new_n806), .B1(new_n780), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n783), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n321), .B1(new_n809), .B2(G329), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n323), .B2(new_n776), .ZN(new_n811));
  INV_X1    g0611(.A(new_n795), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n808), .B(new_n811), .C1(G303), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n802), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n770), .A2(G322), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n791), .B2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT104), .Z(new_n819));
  OAI21_X1  g0619(.A(new_n805), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT105), .ZN(new_n821));
  INV_X1    g0621(.A(new_n764), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n820), .B2(KEYINPUT105), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n767), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n763), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n688), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n751), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  AND2_X1   g0628(.A1(new_n656), .A2(new_n696), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n675), .B1(new_n720), .B2(KEYINPUT26), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n703), .A2(new_n679), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n475), .A2(new_n667), .A3(new_n360), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n468), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n653), .A2(new_n685), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n655), .B1(new_n650), .B2(new_n696), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n653), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n834), .B1(new_n726), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n742), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n752), .B1(new_n838), .B2(new_n742), .ZN(new_n841));
  INV_X1    g0641(.A(new_n837), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n761), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G107), .A2(new_n812), .B1(new_n809), .B2(G311), .ZN(new_n844));
  XNOR2_X1  g0644(.A(KEYINPUT106), .B(G283), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G303), .A2(new_n803), .B1(new_n792), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n773), .ZN(new_n848));
  INV_X1    g0648(.A(new_n780), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n277), .A2(new_n848), .B1(new_n849), .B2(G87), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n321), .B(new_n777), .C1(G294), .C2(new_n770), .ZN(new_n851));
  AND4_X1   g0651(.A1(new_n844), .A2(new_n847), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n776), .A2(new_n201), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G50), .A2(new_n812), .B1(new_n809), .B2(G132), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n321), .C1(new_n202), .C2(new_n780), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n770), .A2(G143), .B1(G159), .B2(new_n848), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n802), .B2(new_n857), .C1(new_n622), .C2(new_n791), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n853), .B(new_n855), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n852), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n822), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n764), .A2(new_n761), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n750), .B(new_n864), .C1(new_n591), .C2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n840), .A2(new_n841), .B1(new_n843), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(G384));
  INV_X1    g0668(.A(new_n389), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n871));
  INV_X1    g0671(.A(G116), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n228), .A2(new_n207), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OAI211_X1 g0675(.A(new_n715), .B(new_n646), .C1(new_n201), .C2(new_n202), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n593), .A2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n206), .B(G13), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n496), .B(new_n281), .C1(new_n880), .C2(KEYINPUT16), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n683), .B1(new_n881), .B2(new_n511), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n662), .B2(new_n532), .ZN(new_n883));
  INV_X1    g0683(.A(new_n530), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n884), .A2(new_n683), .B1(new_n881), .B2(new_n511), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n548), .A2(new_n549), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n557), .A2(new_n683), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT37), .B1(new_n516), .B2(new_n530), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n548), .A4(new_n549), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n883), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n887), .B2(new_n891), .ZN(new_n895));
  INV_X1    g0695(.A(new_n882), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n562), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT107), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n883), .A2(new_n899), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n893), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n601), .A2(new_n685), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n903), .B1(new_n605), .B2(new_n604), .C1(new_n582), .C2(new_n601), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n602), .B2(new_n606), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n835), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n834), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n683), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n901), .A2(new_n909), .B1(new_n659), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT108), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n888), .B1(new_n662), .B2(new_n532), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n531), .A2(new_n546), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT37), .B1(new_n915), .B2(new_n888), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n891), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n913), .B(new_n897), .C1(new_n918), .C2(KEYINPUT38), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n901), .B2(new_n913), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n602), .A2(new_n685), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n659), .A2(new_n910), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n892), .B1(new_n562), .B2(new_n896), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n894), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n883), .A2(new_n899), .A3(new_n895), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n899), .B1(new_n883), .B2(new_n895), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n928), .B2(new_n908), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n912), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n666), .B(new_n725), .C1(new_n726), .C2(KEYINPUT29), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n665), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n932), .B(new_n934), .Z(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n837), .B1(new_n904), .B2(new_n905), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n728), .B2(new_n740), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n901), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n897), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n914), .B2(new_n917), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n938), .B(KEYINPUT40), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n666), .A2(new_n741), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(G330), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n935), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n206), .B2(new_n748), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n935), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n879), .B1(new_n950), .B2(new_n951), .ZN(G367));
  NAND2_X1  g0752(.A1(new_n674), .A2(new_n685), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT112), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n473), .A2(new_n685), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n475), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(new_n702), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n958), .A2(KEYINPUT42), .B1(new_n674), .B2(new_n696), .ZN(new_n959));
  INV_X1    g0759(.A(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n705), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n452), .A2(new_n458), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n685), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n667), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n468), .C2(new_n964), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n959), .A2(new_n962), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT110), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n970), .ZN(new_n972));
  XNOR2_X1  g0772(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT113), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n975), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n969), .A2(new_n975), .A3(new_n974), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n699), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n979), .A2(new_n981), .B1(new_n982), .B2(new_n960), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n977), .A2(new_n978), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n960), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n984), .A2(new_n985), .A3(new_n980), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n706), .A2(new_n708), .A3(new_n957), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT44), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n957), .B1(new_n706), .B2(new_n708), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n982), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n702), .B1(new_n698), .B2(new_n701), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n693), .B(new_n994), .Z(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(new_n699), .A3(new_n991), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n743), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n743), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n712), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n749), .A2(G1), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n987), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n968), .A2(new_n825), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n765), .B1(new_n210), .B2(new_n425), .C1(new_n757), .C2(new_n238), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n752), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G143), .A2(new_n803), .B1(new_n792), .B2(G159), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n776), .A2(new_n202), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n253), .B(new_n1009), .C1(G150), .C2(new_n770), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G58), .A2(new_n812), .B1(new_n809), .B2(G137), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G50), .A2(new_n848), .B1(new_n849), .B2(new_n646), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n323), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G311), .A2(new_n803), .B1(new_n792), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n780), .A2(new_n283), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n795), .A2(new_n1017), .B1(new_n783), .B2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(new_n848), .C2(new_n846), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n776), .A2(new_n341), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n321), .B(new_n1021), .C1(G303), .C2(new_n770), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1015), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT46), .B1(new_n812), .B2(new_n277), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT114), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n1013), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1007), .B1(new_n1027), .B2(new_n764), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1005), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1004), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G387));
  NOR2_X1   g0832(.A1(new_n995), .A2(new_n743), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n712), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n995), .B2(new_n743), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1035), .B2(KEYINPUT117), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT117), .B2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n995), .A2(new_n1002), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n753), .A2(new_n714), .B1(G107), .B2(new_n210), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n235), .A2(new_n264), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n714), .B(new_n264), .C1(new_n202), .C2(new_n591), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n1042));
  NOR3_X1   g0842(.A1(new_n1042), .A2(G50), .A3(new_n507), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(G50), .B2(new_n507), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n757), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n752), .B1(new_n1047), .B2(new_n766), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n771), .A2(new_n593), .B1(new_n215), .B2(new_n795), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n773), .A2(new_n202), .B1(new_n783), .B2(new_n622), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n253), .A4(new_n1016), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n792), .A2(new_n624), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n776), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n427), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n803), .A2(G159), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n321), .B1(new_n809), .B2(G326), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT116), .B(G322), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n803), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n770), .A2(G317), .B1(G303), .B2(new_n848), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n806), .C2(new_n791), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1053), .A2(new_n846), .B1(new_n1014), .B2(new_n812), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1057), .B1(new_n278), .B2(new_n780), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1048), .B1(new_n1070), .B2(new_n764), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n698), .B2(new_n825), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1037), .A2(new_n1038), .A3(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n995), .A2(new_n743), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n996), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n699), .B1(new_n989), .B2(new_n991), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n997), .A3(new_n712), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n756), .A2(new_n245), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n765), .C1(new_n283), .C2(new_n210), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n321), .B(new_n781), .C1(new_n277), .C2(new_n1053), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n792), .A2(G303), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n848), .A2(G294), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n812), .A2(new_n846), .B1(new_n809), .B2(new_n1058), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n803), .A2(G317), .B1(G311), .B2(new_n770), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1053), .A2(G77), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n321), .C1(new_n442), .C2(new_n780), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G68), .A2(new_n812), .B1(new_n809), .B2(G143), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n507), .B2(new_n773), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(G50), .C2(new_n792), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n784), .A2(new_n771), .B1(new_n802), .B2(new_n622), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1088), .A2(new_n1089), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n752), .B(new_n1080), .C1(new_n1097), .C2(new_n822), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n957), .B2(new_n763), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n1002), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1078), .A2(new_n1101), .ZN(G390));
  OAI21_X1  g0902(.A(new_n897), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n921), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n836), .A2(new_n653), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n696), .B(new_n1105), .C1(new_n722), .C2(new_n724), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1106), .A2(new_n907), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1104), .C1(new_n1107), .C2(new_n906), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT119), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n835), .B1(new_n676), .B2(new_n829), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1104), .C1(new_n1110), .C2(new_n906), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT119), .B1(new_n908), .B2(new_n921), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1108), .B1(new_n920), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(G330), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n728), .B2(new_n740), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n906), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n837), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1108), .C1(new_n920), .C2(new_n1113), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1002), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT120), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1116), .A2(new_n666), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n933), .A2(new_n665), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n834), .A2(new_n907), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1117), .B1(new_n1116), .B2(new_n837), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1119), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1129), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n1118), .A3(new_n1107), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1125), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1120), .A2(new_n1121), .A3(new_n1133), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n712), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n865), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n752), .B1(new_n624), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n803), .A2(G128), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n792), .A2(G137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n770), .A2(G132), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n848), .A2(new_n1144), .B1(new_n809), .B2(G125), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n622), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1053), .A2(G159), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n253), .B1(new_n849), .B2(G50), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT53), .B1(new_n795), .B2(new_n622), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n770), .A2(G116), .B1(G294), .B2(new_n809), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G97), .A2(new_n848), .B1(new_n849), .B2(G68), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n796), .A2(new_n321), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n1090), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n802), .A2(new_n807), .B1(new_n791), .B2(new_n341), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1146), .A2(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1139), .B1(new_n1157), .B2(new_n764), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n920), .B2(new_n762), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1124), .A2(new_n1137), .A3(new_n1159), .ZN(G378));
  OAI21_X1  g0960(.A(new_n752), .B1(G50), .B2(new_n1138), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n634), .A2(new_n639), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n630), .A2(new_n683), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(new_n762), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n792), .A2(G97), .B1(new_n427), .B2(new_n848), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n872), .B2(new_n802), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n321), .A2(G41), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n201), .B2(new_n780), .C1(new_n771), .C2(new_n341), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n795), .A2(new_n215), .B1(new_n783), .B2(new_n807), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1174), .A2(new_n1009), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT58), .Z(new_n1179));
  OAI21_X1  g0979(.A(new_n593), .B1(G33), .B2(G41), .ZN(new_n1180));
  INV_X1    g0980(.A(G132), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n791), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n812), .A2(new_n1144), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT121), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n770), .A2(G128), .B1(G137), .B2(new_n848), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n622), .C2(new_n776), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1182), .B(new_n1186), .C1(G125), .C2(new_n803), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT122), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n809), .A2(G124), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n849), .C2(G159), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1179), .B1(new_n1175), .B2(new_n1180), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT123), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n822), .B1(new_n1194), .B2(KEYINPUT123), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1161), .B(new_n1172), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n940), .A2(new_n1171), .A3(G330), .A4(new_n943), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT40), .B1(new_n928), .B2(new_n938), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n943), .A2(G330), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n932), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n921), .A2(new_n920), .B1(new_n929), .B2(new_n930), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1205), .A2(new_n912), .A3(new_n1198), .A4(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1197), .B1(new_n1207), .B2(new_n1002), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1003), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT124), .B1(new_n1211), .B2(new_n1197), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1127), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1136), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1034), .B1(new_n1219), .B2(new_n1215), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT125), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(KEYINPUT125), .B(new_n1034), .C1(new_n1219), .C2(new_n1215), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1213), .B1(new_n1222), .B2(new_n1223), .ZN(G375));
  AND2_X1   g1024(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1127), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1000), .A3(new_n1134), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n750), .B1(new_n202), .B2(new_n865), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT126), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n803), .A2(G294), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1230), .B(new_n1054), .C1(new_n278), .C2(new_n791), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n770), .A2(G283), .B1(G303), .B2(new_n809), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n321), .B1(new_n848), .B2(G107), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n812), .A2(G97), .B1(new_n849), .B2(G77), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n770), .A2(G137), .B1(G159), .B2(new_n812), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G150), .A2(new_n848), .B1(new_n809), .B2(G128), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1053), .A2(G50), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n253), .B1(new_n849), .B2(G58), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n802), .A2(new_n1181), .B1(new_n791), .B2(new_n1143), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1231), .A2(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1229), .B1(new_n764), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1117), .B2(new_n762), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1225), .B2(new_n1003), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1227), .A2(new_n1246), .ZN(G381));
  NOR3_X1   g1047(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n867), .A3(new_n1249), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G387), .A2(G378), .A3(G375), .A4(new_n1250), .ZN(G407));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n684), .A2(G213), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G375), .C2(new_n1255), .ZN(G409));
  OAI211_X1 g1056(.A(G378), .B(new_n1213), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT127), .B1(new_n1216), .B2(new_n999), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1215), .A2(new_n1207), .A3(new_n1259), .A4(new_n1000), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1208), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1252), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1253), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1226), .B1(new_n1133), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1225), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n712), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1246), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n867), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(G384), .A3(new_n1246), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G2897), .A3(new_n1254), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(G2897), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1264), .B2(new_n1272), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(new_n827), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n983), .A2(new_n986), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n999), .B1(new_n997), .B2(new_n743), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1002), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G390), .B1(new_n1284), .B2(new_n1029), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1029), .A3(G390), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1287), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(G396), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(new_n1285), .A3(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1254), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1272), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1278), .A2(new_n1280), .A3(new_n1292), .A4(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1293), .A2(new_n1297), .A3(new_n1294), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1293), .B2(new_n1276), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1296), .B1(new_n1302), .B2(new_n1292), .ZN(G405));
  OR2_X1    g1103(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1252), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1257), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1294), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1272), .A3(new_n1257), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1304), .B(new_n1309), .ZN(G402));
endmodule


