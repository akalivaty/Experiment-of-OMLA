//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G244), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n219), .A2(G77), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  NAND2_X1  g0037(.A1(G68), .A2(G77), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n203), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G222), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n252), .B(new_n254), .C1(new_n202), .C2(new_n253), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT68), .B(G45), .Z(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G41), .A2(G45), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G1), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n207), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n256), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g0068(.A(KEYINPUT69), .B(G226), .Z(new_n269));
  AOI21_X1  g0069(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G200), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT75), .Z(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n216), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n207), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G50), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  INV_X1    g0081(.A(G58), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(KEYINPUT8), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT8), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT71), .A3(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n208), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n279), .A2(new_n282), .A3(new_n201), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n291), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n276), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n280), .B(new_n294), .C1(new_n279), .C2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n257), .A2(G190), .A3(new_n270), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n273), .A2(new_n301), .A3(KEYINPUT10), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n273), .B2(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n284), .A2(G58), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n286), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n289), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n305), .B1(new_n311), .B2(new_n276), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n310), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT73), .A3(new_n275), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n296), .A2(new_n202), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n278), .B2(new_n202), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n253), .A2(G232), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n322), .C1(new_n323), .C2(new_n253), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n256), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n263), .B1(new_n219), .B2(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT72), .B(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n319), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n317), .B1(new_n312), .B2(new_n314), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n327), .A2(G200), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(KEYINPUT74), .B1(G190), .B2(new_n328), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n297), .B1(new_n271), .B2(new_n331), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n257), .A2(new_n329), .A3(new_n270), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n304), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G41), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G1), .A3(G13), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n251), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n261), .A2(new_n262), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n259), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n266), .A2(new_n267), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G238), .A3(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n263), .B1(G238), .B2(new_n268), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n253), .A2(G226), .A3(new_n320), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n349), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n256), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n356), .A2(new_n363), .A3(G179), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT76), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n357), .A2(new_n361), .A3(KEYINPUT76), .A4(new_n362), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(G169), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(KEYINPUT14), .A3(G169), .A4(new_n368), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n365), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n292), .A2(G50), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n375), .B1(new_n208), .B2(G68), .C1(new_n202), .C2(new_n288), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n275), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n276), .A2(G68), .A3(new_n277), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n296), .A2(new_n201), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n367), .A2(G200), .A3(new_n368), .ZN(new_n386));
  INV_X1    g0186(.A(new_n384), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n356), .A2(new_n363), .A3(G190), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT80), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n249), .A2(new_n208), .A3(new_n250), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n249), .A2(new_n394), .A3(new_n208), .A4(new_n250), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(G68), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(G58), .B(G68), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT78), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n396), .A2(new_n402), .A3(KEYINPUT16), .A4(new_n398), .ZN(new_n403));
  AOI211_X1 g0203(.A(new_n276), .B(new_n399), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n287), .A2(new_n277), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT79), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT79), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n287), .A2(new_n407), .A3(new_n277), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n295), .A2(new_n216), .A3(new_n274), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n287), .A2(new_n295), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n391), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n401), .A2(new_n403), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n399), .A2(new_n276), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  OR2_X1    g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G226), .B2(new_n320), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT3), .A2(G33), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT3), .A2(G33), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G87), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n419), .A2(new_n422), .B1(new_n248), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n263), .B1(new_n424), .B2(new_n256), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n268), .A2(G232), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n331), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n329), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n413), .A2(new_n417), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n413), .A2(new_n434), .A3(new_n417), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n414), .A2(new_n415), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n424), .A2(new_n256), .ZN(new_n437));
  AND4_X1   g0237(.A1(G190), .A2(new_n437), .A3(new_n426), .A4(new_n352), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n425), .B2(new_n426), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n412), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n441), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n433), .A2(new_n435), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n345), .A2(new_n390), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G250), .B(new_n320), .C1(new_n420), .C2(new_n421), .ZN(new_n450));
  OAI211_X1 g0250(.A(G257), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G294), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n256), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n455), .A2(new_n347), .A3(G274), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n216), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n455), .A2(new_n457), .B1(new_n459), .B2(new_n346), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G264), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G169), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT87), .ZN(new_n466));
  INV_X1    g0266(.A(G179), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n453), .A2(new_n256), .B1(new_n460), .B2(G264), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT87), .A3(G179), .A4(new_n458), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(KEYINPUT86), .A3(G169), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n468), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n208), .B(G87), .C1(new_n420), .C2(new_n421), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G20), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n208), .B2(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n323), .A2(KEYINPUT23), .A3(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n474), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n275), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT25), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n295), .B2(G107), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n295), .A2(new_n485), .A3(G107), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n207), .A2(G33), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n295), .A2(new_n489), .A3(new_n216), .A4(new_n274), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n487), .A2(new_n488), .B1(new_n323), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT88), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n472), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  INV_X1    g0297(.A(new_n462), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G190), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n462), .A2(G200), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n484), .A2(new_n499), .A3(new_n492), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(G97), .B(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n323), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n393), .A2(G107), .A3(new_n395), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n276), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n296), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n490), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n457), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n347), .ZN(new_n519));
  INV_X1    g0319(.A(G257), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n458), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n320), .C1(new_n420), .C2(new_n421), .ZN(new_n522));
  NOR2_X1   g0322(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n523), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n253), .A2(G244), .A3(new_n320), .A4(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n527));
  AOI22_X1  g0327(.A1(KEYINPUT81), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n521), .B1(new_n529), .B2(new_n256), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT82), .ZN(new_n532));
  OAI21_X1  g0332(.A(G200), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n256), .ZN(new_n534));
  INV_X1    g0334(.A(new_n521), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n534), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n515), .B(new_n531), .C1(new_n533), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n393), .A2(G107), .A3(new_n395), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n292), .A2(G77), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n506), .B1(new_n503), .B2(new_n504), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n208), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n275), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n514), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n538), .A2(new_n331), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n530), .A2(new_n329), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n207), .A2(G45), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G250), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n256), .A2(new_n549), .B1(new_n258), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(G238), .B(new_n320), .C1(new_n420), .C2(new_n421), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n476), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(new_n256), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n439), .ZN(new_n555));
  INV_X1    g0355(.A(G190), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n556), .B(new_n550), .C1(new_n256), .C2(new_n553), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n309), .A2(new_n295), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n490), .A2(new_n423), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n208), .B1(new_n359), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n423), .A2(new_n512), .A3(new_n323), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n208), .B(G68), .C1(new_n420), .C2(new_n421), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n288), .B2(new_n512), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n559), .B(new_n560), .C1(new_n275), .C2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n409), .A2(KEYINPUT83), .A3(new_n309), .A4(new_n489), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  XNOR2_X1  g0370(.A(KEYINPUT15), .B(G87), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n490), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n559), .B1(new_n567), .B2(new_n275), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n554), .B2(new_n329), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n553), .A2(new_n256), .ZN(new_n576));
  INV_X1    g0376(.A(new_n550), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n331), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n558), .A2(new_n568), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n537), .A2(new_n547), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n518), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n258), .B1(new_n459), .B2(new_n346), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n460), .A2(G270), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G264), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n320), .C1(new_n420), .C2(new_n421), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n249), .A2(G303), .A3(new_n250), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n256), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n409), .A2(G116), .A3(new_n489), .ZN(new_n591));
  INV_X1    g0391(.A(G116), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n296), .A2(KEYINPUT84), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n295), .B2(G116), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n274), .A2(new_n216), .B1(G20), .B2(new_n592), .ZN(new_n597));
  NAND2_X1  g0397(.A1(G33), .A2(G283), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n598), .B(new_n208), .C1(G33), .C2(new_n512), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(KEYINPUT20), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT20), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n591), .B(new_n596), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n590), .A2(new_n602), .A3(KEYINPUT21), .A4(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n331), .B1(new_n584), .B2(new_n589), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT85), .A3(KEYINPUT21), .A4(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n602), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n584), .A2(G179), .A3(new_n589), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n609), .A2(new_n610), .B1(new_n602), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n602), .B1(new_n590), .B2(G200), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n556), .B2(new_n590), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n608), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n581), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n502), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n449), .A2(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n573), .A2(new_n574), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n554), .A2(new_n329), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n579), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n608), .A2(new_n612), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n494), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n537), .A2(new_n501), .A3(new_n580), .A4(new_n547), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n511), .A2(new_n514), .B1(new_n530), .B2(G169), .ZN(new_n629));
  INV_X1    g0429(.A(new_n546), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n580), .A3(KEYINPUT26), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT26), .B1(new_n631), .B2(new_n580), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(KEYINPUT89), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n578), .A2(G200), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n554), .A2(G190), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n568), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n545), .A2(new_n546), .A3(new_n621), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n638), .A2(KEYINPUT89), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n628), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n449), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n431), .B(new_n645), .C1(new_n404), .C2(new_n412), .ZN(new_n646));
  INV_X1    g0446(.A(new_n645), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n416), .B2(new_n430), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n374), .A2(new_n384), .B1(new_n389), .B2(new_n333), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n445), .A2(new_n446), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n343), .B1(new_n653), .B2(new_n304), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n644), .A2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n656));
  OAI21_X1  g0456(.A(G213), .B1(new_n656), .B2(KEYINPUT27), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(KEYINPUT27), .B2(new_n656), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT91), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n623), .A2(new_n602), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT92), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n608), .A2(new_n612), .A3(new_n614), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n663), .A2(new_n602), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n664), .B(KEYINPUT92), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n502), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n493), .A2(new_n663), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n468), .A2(new_n470), .ZN(new_n675));
  AOI211_X1 g0475(.A(new_n464), .B(new_n331), .C1(new_n469), .C2(new_n458), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT86), .B1(new_n462), .B2(G169), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n675), .A2(new_n678), .B1(new_n484), .B2(new_n492), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n663), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n671), .A2(KEYINPUT93), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n663), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n624), .A2(new_n663), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n672), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n563), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n214), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n611), .A2(new_n469), .A3(new_n530), .A4(new_n554), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n590), .A2(new_n578), .A3(new_n329), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n538), .A2(new_n462), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n687), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n472), .A2(new_n496), .A3(new_n493), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n496), .B1(new_n472), .B2(new_n493), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n537), .A2(new_n547), .A3(new_n580), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n666), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n710), .A2(new_n501), .A3(new_n712), .A4(new_n687), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n707), .B1(new_n713), .B2(KEYINPUT31), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n705), .B1(new_n704), .B2(KEYINPUT94), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n715), .B(new_n687), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n638), .A2(new_n639), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n633), .A3(KEYINPUT95), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n638), .A2(KEYINPUT95), .A3(new_n639), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n621), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n495), .A2(new_n497), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n627), .B1(new_n727), .B2(new_n623), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n663), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n663), .B1(new_n628), .B2(new_n642), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n721), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n698), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G1), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n693), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n671), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n669), .A2(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n669), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n211), .A2(new_n253), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n211), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n242), .A2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n211), .A2(new_n422), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n215), .B2(new_n261), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n216), .B1(G20), .B2(new_n331), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  OAI21_X1  g0560(.A(new_n742), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n208), .A2(new_n556), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n439), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n208), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G303), .A2(new_n765), .B1(new_n769), .B2(G329), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n766), .A2(new_n763), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n770), .B(new_n422), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n208), .B1(new_n767), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G294), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n762), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n329), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n766), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n329), .A2(new_n779), .A3(new_n439), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G322), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n777), .A2(new_n329), .A3(new_n439), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n329), .A2(new_n779), .A3(G200), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G326), .A2(new_n783), .B1(new_n784), .B2(G311), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n776), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n774), .A2(new_n512), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n780), .B2(G68), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT99), .Z(new_n789));
  NAND2_X1  g0589(.A1(new_n765), .A2(G87), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n253), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT98), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(KEYINPUT98), .B1(G77), .B2(new_n784), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n769), .A2(KEYINPUT32), .A3(G159), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n768), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n772), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n795), .A2(new_n798), .B1(G107), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G50), .A2(new_n783), .B1(new_n778), .B2(G58), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n793), .A2(new_n794), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n786), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n761), .B1(new_n758), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n743), .A2(new_n745), .B1(new_n750), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n758), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n747), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n742), .B1(G77), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT101), .B(G143), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n778), .A2(new_n811), .B1(new_n784), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  INV_X1    g0613(.A(new_n783), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  INV_X1    g0615(.A(new_n780), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n812), .B1(new_n813), .B2(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n253), .B1(new_n764), .B2(new_n279), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n799), .A2(G68), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n768), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(G58), .C2(new_n775), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G116), .A2(new_n784), .B1(new_n780), .B2(G283), .ZN(new_n827));
  INV_X1    g0627(.A(G303), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n814), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT100), .Z(new_n830));
  NOR2_X1   g0630(.A1(new_n772), .A2(new_n423), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G311), .B2(new_n769), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(new_n422), .C1(new_n323), .C2(new_n764), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n787), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  INV_X1    g0635(.A(new_n778), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n826), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n807), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n809), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n337), .A2(new_n339), .ZN(new_n843));
  INV_X1    g0643(.A(new_n333), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n319), .A2(new_n663), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n319), .A2(new_n330), .A3(new_n663), .A4(new_n332), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n747), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n721), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n340), .A2(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n732), .B(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n742), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n853), .A2(new_n856), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n739), .A2(new_n207), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n663), .A2(new_n384), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n389), .B(new_n862), .C1(new_n373), .C2(new_n387), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n373), .A2(new_n862), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n854), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n714), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT80), .B1(new_n436), .B2(new_n442), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n391), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(new_n661), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n443), .B1(new_n416), .B2(new_n430), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n661), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n413), .A2(new_n417), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n432), .A2(new_n875), .A3(new_n876), .A4(new_n443), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n871), .B1(new_n649), .B2(new_n652), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n436), .B2(new_n442), .ZN(new_n884));
  AOI211_X1 g0684(.A(KEYINPUT104), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n431), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n443), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n877), .ZN(new_n890));
  INV_X1    g0690(.A(new_n886), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n448), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n868), .A2(KEYINPUT106), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n652), .B1(KEYINPUT18), .B2(new_n432), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n886), .B1(new_n896), .B2(new_n435), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n443), .A2(new_n876), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n869), .A2(new_n870), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n431), .ZN(new_n900));
  AOI22_X1  g0700(.A1(KEYINPUT37), .A2(new_n888), .B1(new_n900), .B2(new_n875), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n881), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n902), .A2(new_n895), .A3(new_n893), .ZN(new_n903));
  NAND2_X1  g0703(.A1(KEYINPUT106), .A2(KEYINPUT40), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n865), .B(new_n904), .C1(new_n714), .C2(new_n867), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n894), .A2(new_n895), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n449), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n714), .A2(new_n867), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n715), .B1(new_n617), .B2(new_n687), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n866), .B1(new_n911), .B2(new_n707), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n449), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n913), .A3(G330), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n374), .A2(new_n384), .A3(new_n687), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n878), .B2(new_n879), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n889), .A2(new_n877), .B1(new_n448), .B2(new_n891), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(KEYINPUT38), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n915), .B(new_n918), .C1(new_n921), .C2(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n902), .A2(new_n893), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n863), .A2(new_n864), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT89), .B1(new_n638), .B2(new_n639), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n722), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n640), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n679), .A2(new_n623), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n621), .B1(new_n928), .B2(new_n626), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n687), .B(new_n851), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n844), .A2(new_n663), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n924), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n923), .A2(new_n933), .B1(new_n649), .B2(new_n661), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n449), .B1(new_n734), .B2(new_n731), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n654), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n861), .B1(new_n914), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n914), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(G116), .A4(new_n217), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT36), .ZN(new_n944));
  OAI21_X1  g0744(.A(G77), .B1(new_n282), .B2(new_n201), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n945), .A2(new_n214), .B1(G50), .B2(new_n201), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n737), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n944), .A3(new_n947), .ZN(G367));
  INV_X1    g0748(.A(new_n760), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n211), .B2(new_n571), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n236), .A2(new_n755), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n742), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G317), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n422), .B1(new_n768), .B2(new_n953), .C1(new_n512), .C2(new_n772), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n764), .B2(new_n592), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n323), .C2(new_n774), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n954), .B(new_n958), .C1(G294), .C2(new_n780), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G303), .A2(new_n778), .B1(new_n783), .B2(G311), .ZN(new_n960));
  INV_X1    g0760(.A(new_n784), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n960), .C1(new_n771), .C2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G58), .A2(new_n765), .B1(new_n769), .B2(G137), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n772), .A2(new_n202), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n422), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n775), .A2(G68), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n783), .A2(new_n811), .B1(new_n784), .B2(G50), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n815), .B2(new_n836), .C1(new_n797), .C2(new_n816), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n952), .B1(new_n971), .B2(new_n758), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n687), .A2(new_n568), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT107), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(new_n622), .ZN(new_n975));
  INV_X1    g0775(.A(new_n580), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n972), .B1(new_n979), .B2(new_n749), .ZN(new_n980));
  INV_X1    g0780(.A(new_n686), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n537), .B(new_n547), .C1(new_n515), .C2(new_n687), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n631), .A2(new_n663), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n690), .A2(new_n688), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT45), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n690), .A2(new_n688), .ZN(new_n987));
  INV_X1    g0787(.A(new_n984), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT44), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n987), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n981), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n686), .B(new_n986), .C1(new_n989), .C2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT109), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n681), .A2(new_n994), .A3(new_n689), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n681), .B2(new_n689), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n690), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n671), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n995), .A2(new_n670), .A3(new_n690), .A4(new_n996), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n992), .A2(new_n993), .A3(new_n735), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n735), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n693), .B(KEYINPUT41), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n741), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n672), .A2(new_n689), .A3(new_n984), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n727), .A2(new_n537), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n687), .B1(new_n1010), .B2(new_n631), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT108), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n978), .B(KEYINPUT43), .Z(new_n1017));
  OAI22_X1  g0817(.A1(new_n1014), .A2(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n981), .A2(new_n984), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n980), .B1(new_n1005), .B2(new_n1022), .ZN(G387));
  AOI21_X1  g0823(.A(new_n694), .B1(new_n1000), .B2(new_n735), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n735), .B2(new_n1000), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n233), .A2(new_n261), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(new_n755), .B1(new_n695), .B2(new_n751), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n307), .A2(new_n279), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT50), .Z(new_n1029));
  NAND4_X1  g0829(.A1(new_n1029), .A2(new_n456), .A3(new_n238), .A4(new_n695), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1027), .A2(new_n1030), .B1(new_n323), .B2(new_n692), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n742), .B1(new_n1031), .B2(new_n760), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G159), .A2(new_n783), .B1(new_n784), .B2(G68), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G50), .A2(new_n778), .B1(new_n780), .B2(new_n287), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n764), .A2(new_n202), .B1(new_n768), .B2(new_n815), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n253), .B1(new_n772), .B2(new_n512), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n774), .A2(new_n571), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n253), .B1(new_n769), .B2(G326), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G322), .A2(new_n783), .B1(new_n780), .B2(G311), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT111), .Z(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n828), .B2(new_n961), .C1(new_n953), .C2(new_n836), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n765), .A2(G294), .B1(new_n775), .B2(G283), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1040), .B1(new_n592), .B2(new_n772), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1032), .B1(new_n1052), .B2(new_n758), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n681), .B2(new_n749), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1025), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1000), .A2(new_n741), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT110), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1055), .A2(new_n1057), .ZN(G393));
  NAND3_X1  g0858(.A1(new_n992), .A2(new_n993), .A3(new_n741), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n988), .A2(new_n748), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT112), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n742), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n778), .B1(new_n783), .B2(G317), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  AOI22_X1  g0864(.A1(G283), .A2(new_n765), .B1(new_n769), .B2(G322), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n422), .C1(new_n323), .C2(new_n772), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G116), .B2(new_n775), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G294), .A2(new_n784), .B1(new_n780), .B2(G303), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n783), .B1(new_n778), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  OAI22_X1  g0871(.A1(new_n810), .A2(new_n768), .B1(new_n764), .B2(new_n201), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n774), .A2(new_n202), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1072), .A2(new_n831), .A3(new_n1073), .A4(new_n422), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G50), .A2(new_n780), .B1(new_n784), .B2(new_n307), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n807), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n245), .A2(new_n211), .A3(new_n422), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n760), .B1(G97), .B2(new_n692), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1062), .B(new_n1077), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1061), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1001), .A2(new_n693), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n992), .A2(new_n993), .B1(new_n735), .B2(new_n1000), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1059), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(G390));
  OAI21_X1  g0884(.A(KEYINPUT113), .B1(new_n933), .B2(new_n918), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n916), .B(KEYINPUT105), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n931), .B1(new_n732), .B2(new_n851), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1087), .C1(new_n1088), .C2(new_n924), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n915), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT39), .B1(new_n882), .B2(new_n893), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1085), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n882), .A2(new_n893), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n931), .B1(new_n729), .B2(new_n851), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1087), .C1(new_n1094), .C2(new_n924), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n912), .A2(KEYINPUT114), .A3(G330), .A4(new_n865), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n865), .B(G330), .C1(new_n714), .C2(new_n867), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n865), .B(G330), .C1(new_n714), .C2(new_n718), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1092), .A2(new_n1103), .A3(new_n1095), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n741), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT115), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1102), .A2(new_n1108), .A3(new_n741), .A4(new_n1104), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n909), .A2(new_n720), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n449), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n936), .A3(new_n654), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n851), .C1(new_n714), .C2(new_n718), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n924), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1097), .A2(new_n1100), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1088), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n912), .A2(G330), .A3(new_n851), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n924), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1113), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1105), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1102), .A2(new_n1123), .A3(new_n1104), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n693), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n746), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n742), .B1(new_n287), .B2(new_n808), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n813), .A2(new_n816), .B1(new_n961), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G128), .B2(new_n783), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT53), .B1(new_n764), .B2(new_n815), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G159), .B2(new_n775), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n422), .B1(new_n769), .B2(G125), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n279), .B2(new_n772), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G132), .B2(new_n778), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G97), .A2(new_n784), .B1(new_n780), .B2(G107), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n771), .B2(new_n814), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT116), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n769), .A2(G294), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n790), .A2(new_n822), .A3(new_n1143), .A4(new_n422), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n1073), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n592), .B2(new_n836), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1129), .B1(new_n1147), .B2(new_n758), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1128), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1110), .A2(new_n1127), .A3(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n304), .A2(new_n344), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n297), .A2(new_n661), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n935), .A2(new_n906), .A3(G330), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n935), .B1(G330), .B2(new_n906), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n906), .A2(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n922), .A3(new_n934), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1160), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1161), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1106), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n746), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n742), .B1(G50), .B2(new_n808), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n764), .A2(new_n1130), .B1(new_n774), .B2(new_n815), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G128), .A2(new_n778), .B1(new_n784), .B2(G137), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n823), .B2(new_n816), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G125), .C2(new_n783), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT59), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n799), .A2(G159), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G41), .B(new_n253), .C1(new_n765), .C2(G77), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n769), .A2(G283), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n799), .A2(G58), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n966), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n323), .A2(new_n836), .B1(new_n816), .B2(new_n512), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n592), .A2(new_n814), .B1(new_n961), .B2(new_n571), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n279), .B1(new_n420), .B2(G41), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1181), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1171), .B1(new_n1193), .B2(new_n758), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1170), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT118), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT118), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1170), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT119), .B1(new_n1169), .B2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1162), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1167), .B1(new_n1166), .B2(new_n1161), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n741), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1199), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT119), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1113), .B(KEYINPUT120), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1164), .A2(new_n1168), .B1(new_n1126), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n693), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1126), .A2(new_n1207), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1200), .B(new_n1206), .C1(new_n1209), .C2(new_n1212), .ZN(G375));
  AOI22_X1  g1013(.A1(new_n1116), .A2(new_n1117), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1113), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1124), .A2(new_n1004), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n924), .A2(new_n746), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n742), .B1(G68), .B2(new_n808), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n764), .A2(new_n512), .B1(new_n768), .B2(new_n828), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1219), .A2(new_n964), .A3(new_n1037), .A4(new_n253), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G107), .A2(new_n784), .B1(new_n780), .B2(G116), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G283), .A2(new_n778), .B1(new_n783), .B2(G294), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n784), .A2(G150), .B1(G50), .B2(new_n775), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  AOI22_X1  g1025(.A1(G159), .A2(new_n765), .B1(new_n769), .B2(G128), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(new_n253), .A3(new_n1184), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1130), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G137), .A2(new_n778), .B1(new_n780), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(new_n823), .C2(new_n814), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1218), .B1(new_n1231), .B2(new_n758), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1217), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1214), .B2(new_n1106), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1216), .A2(new_n1235), .ZN(G381));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  INV_X1    g1037(.A(G384), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OR3_X1    g1039(.A1(new_n1055), .A2(new_n1057), .A3(G396), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1239), .A2(G387), .A3(new_n1240), .A4(G381), .ZN(new_n1241));
  INV_X1    g1041(.A(G378), .ZN(new_n1242));
  INV_X1    g1042(.A(G375), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1242), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(new_n1245), .C2(G343), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(G409));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G387), .B2(new_n1237), .ZN(new_n1249));
  OAI21_X1  g1049(.A(G396), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1240), .A2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G387), .A2(new_n1237), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1003), .B1(new_n1001), .B2(new_n735), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1021), .B(new_n1020), .C1(new_n1253), .C2(new_n741), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G390), .B1(new_n1254), .B2(new_n980), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1249), .A2(new_n1251), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1240), .A2(new_n1250), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(new_n1237), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1254), .A2(new_n980), .A3(G390), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1248), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1206), .A2(new_n1200), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G378), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1210), .A2(new_n1004), .A3(new_n1211), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1265), .A2(new_n1203), .A3(new_n1195), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1266), .A2(new_n1242), .B1(G213), .B2(new_n662), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1124), .A2(new_n693), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT60), .B1(new_n1215), .B2(KEYINPUT123), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1215), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1273), .A2(new_n1238), .A3(new_n1234), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1215), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n693), .B(new_n1124), .C1(new_n1275), .C2(new_n1270), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1276), .B2(new_n1235), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1274), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1238), .B1(new_n1273), .B2(new_n1234), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1276), .A2(G384), .A3(new_n1235), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1264), .A2(new_n1267), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1261), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1283), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1281), .A2(new_n1282), .A3(new_n1278), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n662), .A2(G213), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1265), .A2(new_n1203), .A3(new_n1195), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(G378), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(G378), .B2(G375), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1300), .B2(new_n1286), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1264), .A2(new_n1267), .A3(KEYINPUT63), .A4(new_n1286), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1292), .B1(new_n1303), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1287), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1285), .A2(new_n1310), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1311), .A2(KEYINPUT125), .A3(new_n1306), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1291), .B1(new_n1308), .B2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1314));
  OR3_X1    g1114(.A1(new_n1314), .A2(KEYINPUT126), .A3(KEYINPUT127), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT127), .B1(new_n1314), .B2(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1304), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1261), .A2(new_n1316), .A3(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1245), .A2(new_n1264), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(KEYINPUT126), .B2(new_n1314), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1320), .B(new_n1322), .ZN(G402));
endmodule


