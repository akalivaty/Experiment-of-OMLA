//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n465), .A2(G2104), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G2105), .B1(G101), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g062(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n465), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n471), .A2(G136), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n465), .C1(new_n475), .C2(new_n476), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n464), .A2(new_n501), .A3(G138), .A4(new_n465), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT72), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G88), .B1(new_n515), .B2(G50), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n506), .A2(new_n508), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(KEYINPUT73), .A3(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n525), .A2(KEYINPUT74), .A3(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT74), .B1(new_n525), .B2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n512), .A2(G51), .A3(G543), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT75), .B(G89), .Z(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n509), .A2(new_n512), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n514), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n542), .A2(new_n549), .B1(new_n514), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n520), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n513), .B2(G91), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n563), .B(G543), .C1(new_n511), .C2(new_n510), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n528), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT77), .B(new_n516), .C1(new_n526), .C2(new_n527), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(G303));
  NAND2_X1  g146(.A1(new_n513), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n515), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n542), .A2(new_n576), .B1(new_n514), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n509), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT78), .Z(new_n581));
  AOI21_X1  g156(.A(new_n540), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n520), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n590), .A3(G651), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT80), .B(G47), .Z(new_n592));
  AOI22_X1  g167(.A1(new_n513), .A2(G85), .B1(new_n515), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n540), .B1(new_n597), .B2(new_n514), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI221_X1 g175(.A(KEYINPUT81), .B1(new_n514), .B2(new_n597), .C1(new_n596), .C2(new_n540), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n542), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT10), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n464), .A2(new_n480), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n484), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n471), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n465), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n623), .A2(new_n624), .A3(new_n631), .ZN(G156));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  OAI21_X1  g211(.A(KEYINPUT14), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n643), .A2(new_n648), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(G14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(new_n653), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n658), .B2(new_n651), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n622), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n630), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT86), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n675), .A2(new_n676), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n678), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n674), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n687), .B1(new_n683), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  OR3_X1    g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n688), .B2(new_n689), .ZN(new_n693));
  AND3_X1   g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n583), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT33), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT33), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1976), .ZN(new_n708));
  INV_X1    g283(.A(G1976), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n700), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n701), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n701), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT89), .B(G1971), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n714), .A2(new_n716), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n711), .A2(new_n712), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n701), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n701), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1986), .Z(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n484), .A2(G119), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT88), .Z(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G131), .B2(new_n471), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(new_n724), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n719), .A2(new_n723), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n711), .A2(new_n717), .A3(new_n718), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(KEYINPUT90), .A3(KEYINPUT34), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n737), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n737), .A2(new_n741), .A3(new_n742), .A4(new_n745), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G129), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G105), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n471), .A2(G141), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT26), .Z(new_n759));
  NAND4_X1  g334(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n724), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n724), .B2(G32), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n754), .B1(new_n724), .B2(new_n629), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n724), .A2(G27), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n724), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G2078), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n701), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n701), .B2(G21), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(G2078), .B2(new_n768), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT24), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(KEYINPUT97), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT97), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n482), .B2(new_n724), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2084), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n766), .A2(new_n769), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G171), .A2(new_n701), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G5), .B2(new_n701), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n724), .A2(G26), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT28), .Z(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n789));
  OAI211_X1 g364(.A(G128), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n471), .B2(G140), .ZN(new_n793));
  OAI211_X1 g368(.A(G140), .B(new_n465), .C1(new_n475), .C2(new_n476), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n791), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n787), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n783), .A2(new_n784), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n701), .A2(G19), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n552), .B2(new_n701), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G1341), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n785), .A2(new_n798), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n781), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n771), .A2(new_n772), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT98), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n724), .A2(G33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n471), .A2(G139), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n465), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT25), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n810), .A2(new_n815), .A3(KEYINPUT96), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT96), .B1(new_n810), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n807), .B1(new_n818), .B2(new_n724), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G2072), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(G2072), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n806), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G4), .A2(G16), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT93), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n606), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1348), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n801), .A2(G1341), .ZN(new_n827));
  NOR2_X1   g402(.A1(G29), .A2(G35), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G162), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2090), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n701), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1956), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n832), .B(new_n836), .C1(new_n831), .C2(new_n830), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n804), .A2(new_n822), .A3(new_n826), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n747), .A2(new_n748), .A3(new_n838), .ZN(G311));
  NAND3_X1  g414(.A1(new_n747), .A2(new_n748), .A3(new_n838), .ZN(G150));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n542), .A2(new_n841), .B1(new_n514), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n509), .A2(G67), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n540), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n845), .B1(new_n520), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G651), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n513), .A2(G93), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n515), .A2(G55), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n853), .A2(KEYINPUT100), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n843), .B2(new_n846), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n856), .B(new_n858), .C1(new_n548), .C2(new_n551), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n552), .A2(new_n847), .A3(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n606), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n848), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n850), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT101), .ZN(G145));
  NAND2_X1  g445(.A1(new_n484), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n465), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G142), .B2(new_n471), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT107), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n732), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n493), .A2(new_n497), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(KEYINPUT103), .B1(new_n500), .B2(new_n502), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n498), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n796), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n500), .A2(new_n502), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n493), .A2(KEYINPUT103), .A3(new_n497), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n789), .A2(new_n790), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n471), .A2(new_n792), .A3(G140), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n884), .A2(new_n892), .A3(new_n761), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n761), .B1(new_n884), .B2(new_n892), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT104), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n796), .B1(new_n881), .B2(new_n883), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n887), .A2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n760), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n884), .A2(new_n892), .A3(new_n761), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n879), .B(new_n818), .C1(new_n895), .C2(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n818), .A2(new_n893), .A3(new_n894), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n818), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT104), .B1(new_n893), .B2(new_n894), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n899), .A2(new_n896), .A3(new_n900), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(new_n879), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n620), .B(KEYINPUT106), .Z(new_n911));
  NOR3_X1   g486(.A1(new_n905), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n903), .B1(new_n909), .B2(new_n879), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n818), .B1(new_n895), .B2(new_n901), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n878), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n911), .B1(new_n905), .B2(new_n910), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n916), .A3(new_n913), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n877), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n629), .B(KEYINPUT102), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(G162), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n482), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n918), .A2(new_n925), .A3(new_n921), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT40), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n919), .A2(new_n877), .A3(new_n920), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n877), .B1(new_n919), .B2(new_n920), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  AND4_X1   g508(.A1(KEYINPUT40), .A2(new_n932), .A3(new_n933), .A4(new_n928), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n929), .A2(new_n934), .ZN(G395));
  XNOR2_X1  g510(.A(new_n615), .B(new_n861), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n602), .A2(G299), .A3(new_n605), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G299), .B1(new_n602), .B2(new_n605), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n602), .A2(new_n605), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n610), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n937), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n936), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n528), .A2(new_n721), .ZN(new_n951));
  OAI211_X1 g526(.A(G290), .B(new_n516), .C1(new_n526), .C2(new_n527), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n583), .B(G288), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n953), .B(new_n954), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT109), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n949), .A2(new_n950), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n946), .A2(new_n948), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n958), .A2(new_n959), .B1(KEYINPUT110), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n957), .ZN(new_n962));
  AND4_X1   g537(.A1(KEYINPUT110), .A2(new_n960), .A3(new_n962), .A4(new_n959), .ZN(new_n963));
  OAI21_X1  g538(.A(G868), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n847), .A2(G868), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G295));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n965), .ZN(G331));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g543(.A1(G301), .A2(G286), .ZN(new_n969));
  NAND2_X1  g544(.A1(G168), .A2(G171), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n861), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n859), .A2(new_n860), .A3(new_n969), .A4(new_n970), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n947), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n941), .B2(new_n944), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n947), .A2(new_n972), .A3(KEYINPUT111), .A4(new_n973), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n955), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n953), .B(new_n954), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n933), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n975), .A2(new_n987), .A3(KEYINPUT41), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT41), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n947), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n974), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n972), .A2(new_n973), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n947), .B1(new_n992), .B2(new_n940), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n955), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n933), .A4(new_n983), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n985), .A2(new_n986), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n983), .A2(new_n933), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n996), .A4(new_n980), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n980), .A2(new_n996), .A3(new_n933), .A4(new_n983), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT113), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n982), .B1(new_n991), .B2(new_n993), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n984), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n998), .B1(new_n1006), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n887), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n473), .A2(G40), .A3(new_n481), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n732), .B(new_n735), .Z(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n760), .B(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n891), .B(G2067), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G290), .A2(G1986), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1012), .A3(KEYINPUT48), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(new_n1011), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1018), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1011), .A2(G1996), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT46), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1011), .B1(new_n761), .B2(new_n1016), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n733), .A2(new_n735), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1030), .A2(new_n1017), .B1(G2067), .B2(new_n796), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1024), .B(new_n1029), .C1(new_n1012), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n887), .A2(new_n1008), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n473), .A2(new_n481), .A3(G40), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n583), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G1981), .B1(new_n578), .B2(new_n582), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n1035), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n709), .A3(new_n703), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1035), .B1(new_n1046), .B2(new_n1037), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(G164), .B2(G1384), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1010), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1971), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n885), .A2(new_n880), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1008), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT50), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n887), .A2(new_n1058), .A3(new_n1008), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1010), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2090), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n569), .A2(G8), .A3(new_n570), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n569), .A2(KEYINPUT55), .A3(G8), .A4(new_n570), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT118), .B(G8), .C1(new_n1054), .C2(new_n1061), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n703), .B2(G1976), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G288), .A2(new_n709), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1035), .A3(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1035), .A2(new_n1073), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(KEYINPUT52), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1045), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(G164), .A2(new_n1049), .A3(G1384), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1009), .A2(new_n1079), .A3(new_n1034), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n772), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1057), .A2(new_n1010), .A3(new_n1059), .ZN(new_n1083));
  INV_X1    g658(.A(G2084), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G168), .A2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1070), .A2(new_n1078), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1047), .B1(new_n1089), .B2(KEYINPUT63), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1055), .A2(new_n1058), .A3(new_n1008), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g667(.A(G2090), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1034), .B1(new_n1033), .B2(KEYINPUT50), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1053), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1067), .B(new_n1068), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1086), .A2(KEYINPUT63), .A3(new_n1087), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1062), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1101), .A2(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1090), .B1(new_n1105), .B2(new_n1077), .ZN(new_n1106));
  OAI221_X1 g681(.A(G168), .B1(new_n1060), .B2(G2084), .C1(new_n1080), .C2(G1966), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(G168), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1111), .A3(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT62), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(G2078), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1080), .A2(new_n1116), .B1(new_n1060), .B2(new_n784), .ZN(new_n1117));
  INV_X1    g692(.A(G2078), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1048), .A2(new_n1010), .A3(new_n1118), .A4(new_n1050), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1115), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1119), .B2(new_n1115), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G171), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1110), .A2(new_n1127), .A3(new_n1112), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1114), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1121), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(G301), .A3(new_n1117), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n1083), .B2(G1961), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1060), .A2(new_n1134), .A3(new_n784), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n1009), .A2(KEYINPUT126), .A3(new_n1034), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n1009), .B2(new_n1034), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1048), .A3(new_n1116), .A4(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1131), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT54), .B(new_n1132), .C1(new_n1140), .C2(G301), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1131), .A2(new_n1136), .A3(G301), .A4(new_n1139), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1142), .A2(KEYINPUT127), .A3(new_n1125), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1142), .B2(KEYINPUT127), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1141), .B(new_n1113), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1956), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1148));
  INV_X1    g723(.A(G91), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1148), .A2(new_n540), .B1(new_n542), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT120), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n560), .A2(G651), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n513), .A2(G91), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1155), .A3(new_n565), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1157));
  NAND4_X1  g732(.A1(new_n1152), .A2(KEYINPUT57), .A3(new_n1154), .A4(new_n565), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT121), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n561), .A2(new_n1160), .A3(KEYINPUT57), .A4(new_n565), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1156), .A2(new_n1157), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT56), .B(G2072), .Z(new_n1163));
  NOR2_X1   g738(.A1(new_n1051), .A2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1147), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1348), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1060), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G2067), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1010), .A2(new_n1008), .A3(new_n1168), .A4(new_n887), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n606), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1162), .B1(new_n1147), .B2(new_n1164), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1165), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n606), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n942), .A4(new_n1169), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1175), .A2(new_n1176), .B1(new_n1177), .B2(new_n1170), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(G1956), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT116), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1091), .B(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1094), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1164), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1181), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT123), .B1(new_n1165), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1178), .B1(new_n1189), .B2(KEYINPUT61), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1186), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n1172), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1048), .A2(new_n1010), .A3(new_n1014), .A4(new_n1050), .ZN(new_n1195));
  XOR2_X1   g770(.A(KEYINPUT58), .B(G1341), .Z(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n552), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT59), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT59), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1193), .A2(new_n1194), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1173), .B1(new_n1190), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1129), .B1(new_n1146), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1077), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1101), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1106), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(G290), .B(G1986), .Z(new_n1211));
  OAI21_X1  g786(.A(new_n1018), .B1(new_n1011), .B2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT114), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1032), .B1(new_n1210), .B2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g789(.A1(G227), .A2(new_n461), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1216), .B1(new_n694), .B2(new_n695), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1217), .B1(new_n656), .B2(new_n659), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n996), .B1(new_n999), .B2(new_n980), .ZN(new_n1219));
  NOR3_X1   g793(.A1(new_n984), .A2(KEYINPUT43), .A3(new_n1004), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n928), .B2(new_n927), .ZN(G308));
  NAND2_X1  g796(.A1(new_n927), .A2(new_n928), .ZN(new_n1223));
  OAI211_X1 g797(.A(new_n1223), .B(new_n1218), .C1(new_n1219), .C2(new_n1220), .ZN(G225));
endmodule


