//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n466), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n466), .A2(new_n468), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT65), .B(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n464), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND2_X1  g069(.A1(new_n479), .A2(G102), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n477), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n475), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n464), .A2(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n467), .A2(G2104), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n498), .B(new_n502), .C1(new_n508), .C2(KEYINPUT4), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n512), .A2(new_n514), .A3(new_n519), .A4(new_n521), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n518), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  INV_X1    g104(.A(new_n523), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  INV_X1    g106(.A(new_n526), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n517), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n523), .A2(new_n541), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n517), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n523), .A2(new_n547), .B1(new_n548), .B2(new_n526), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n561), .A2(new_n517), .B1(new_n562), .B2(new_n526), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n560), .B1(new_n559), .B2(new_n563), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G49), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n523), .A2(new_n569), .B1(new_n570), .B2(new_n526), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g149(.A(KEYINPUT69), .B(G651), .C1(new_n515), .C2(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n512), .A2(new_n514), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n515), .A2(new_n522), .A3(G86), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n519), .A2(new_n521), .A3(G48), .A4(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n512), .A2(new_n514), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(KEYINPUT70), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(KEYINPUT70), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(G651), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT71), .B(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n530), .A2(new_n592), .B1(G85), .B2(new_n532), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n530), .A2(G54), .B1(new_n598), .B2(G651), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n526), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g176(.A(KEYINPUT72), .B(KEYINPUT10), .Z(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT73), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n488), .A2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n490), .A2(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT76), .B(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n506), .A2(new_n507), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n479), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT77), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT78), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  OAI211_X1 g231(.A(KEYINPUT17), .B(new_n653), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n654), .ZN(new_n660));
  OAI221_X1 g235(.A(new_n657), .B1(new_n658), .B2(new_n654), .C1(new_n660), .C2(new_n653), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n653), .A3(new_n656), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(KEYINPUT81), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(KEYINPUT81), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n669), .A2(new_n670), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n676), .A2(new_n681), .A3(new_n672), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G229));
  XNOR2_X1  g265(.A(KEYINPUT35), .B(G1991), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n488), .A2(G119), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n490), .A2(G131), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  NOR2_X1   g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT85), .Z(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT86), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n694), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n704));
  OR2_X1    g279(.A1(G25), .A2(G29), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n692), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n703), .A2(new_n705), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT87), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n711), .A2(new_n691), .A3(new_n706), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n576), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G16), .B2(G23), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT33), .B(G1976), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n714), .A2(G6), .ZN(new_n722));
  INV_X1    g297(.A(G305), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n714), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT32), .B(G1981), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT88), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n717), .A2(new_n721), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n717), .A2(KEYINPUT34), .A3(new_n721), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G290), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G24), .ZN(new_n735));
  INV_X1    g310(.A(G1986), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n713), .A2(new_n732), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT36), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n709), .A2(new_n712), .B1(new_n736), .B2(new_n735), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n741), .A2(new_n742), .A3(new_n732), .A4(new_n737), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G164), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G27), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n702), .A2(G26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n490), .A2(G140), .ZN(new_n751));
  OAI221_X1 g326(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT90), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(G29), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n749), .B(new_n755), .S(KEYINPUT28), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  AND2_X1   g332(.A1(KEYINPUT30), .A2(G28), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT30), .A2(G28), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n702), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(new_n626), .C2(new_n702), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  NOR2_X1   g338(.A1(new_n746), .A2(new_n747), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n714), .A2(KEYINPUT23), .A3(G20), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G20), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G16), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n769), .C1(new_n610), .C2(new_n714), .ZN(new_n770));
  INV_X1    g345(.A(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n714), .A2(G4), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n606), .B2(new_n714), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT89), .B(G1348), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n757), .A2(new_n765), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n702), .A2(G33), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n629), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n464), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT91), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n490), .A2(G139), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT25), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n781), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(new_n702), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G2072), .Z(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G35), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G162), .B2(G29), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT29), .B(G2090), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G21), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G168), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT93), .B(G1966), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n714), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n550), .B2(new_n714), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(G1341), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(G1341), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n797), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G5), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G171), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1961), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n795), .B2(new_n796), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n789), .A2(new_n793), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n777), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n744), .A2(new_n748), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n490), .A2(G141), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n479), .A2(G105), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT26), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n813), .B(new_n815), .C1(new_n488), .C2(G129), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G29), .B2(G32), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT27), .B(G1996), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(KEYINPUT24), .A2(G34), .ZN(new_n824));
  NAND2_X1  g399(.A1(KEYINPUT24), .A2(G34), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n702), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G160), .B2(new_n702), .ZN(new_n827));
  INV_X1    g402(.A(G2084), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n809), .A2(KEYINPUT95), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n744), .A2(new_n808), .A3(new_n829), .A4(new_n748), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n822), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n833), .ZN(G311));
  NAND3_X1  g409(.A1(new_n809), .A2(new_n823), .A3(new_n829), .ZN(G150));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT97), .B(G93), .Z(new_n837));
  OAI22_X1  g412(.A1(new_n523), .A2(new_n836), .B1(new_n526), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n515), .A2(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n517), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n606), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(KEYINPUT98), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n838), .A2(new_n841), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n550), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n550), .A3(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n847), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n845), .B1(new_n859), .B2(G860), .ZN(G145));
  NAND2_X1  g435(.A1(new_n488), .A2(G130), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n490), .A2(G142), .ZN(new_n862));
  OAI221_X1 g437(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n701), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n817), .B(new_n509), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n865), .B(new_n866), .Z(new_n867));
  INV_X1    g442(.A(G160), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n868), .A3(new_n625), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n624), .B2(new_n625), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n493), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(G162), .A3(new_n869), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n874), .A3(new_n786), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n786), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n754), .B(new_n631), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n865), .B(new_n866), .ZN(new_n880));
  INV_X1    g455(.A(new_n877), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n879), .B1(new_n878), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g463(.A(new_n856), .B(new_n615), .Z(new_n889));
  INV_X1    g464(.A(new_n566), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT100), .B1(new_n890), .B2(new_n564), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n565), .A2(new_n892), .A3(new_n566), .ZN(new_n893));
  INV_X1    g468(.A(new_n605), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(G299), .A2(KEYINPUT100), .A3(new_n605), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G290), .A2(G303), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(G290), .A2(G303), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n723), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(G305), .A3(new_n905), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n908), .A2(new_n910), .A3(new_n576), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n576), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n904), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G868), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n849), .A2(G868), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(G295));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n922), .ZN(new_n925));
  AOI211_X1 g500(.A(KEYINPUT102), .B(new_n921), .C1(new_n919), .C2(G868), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  XNOR2_X1  g503(.A(G286), .B(G171), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n854), .A2(new_n928), .A3(new_n855), .A4(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  INV_X1    g506(.A(new_n855), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n550), .B1(new_n848), .B2(new_n851), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n854), .A2(new_n855), .A3(new_n929), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT103), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n901), .A2(new_n902), .A3(new_n930), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n898), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n913), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(new_n913), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n937), .A2(new_n945), .A3(new_n913), .A4(new_n939), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n941), .A2(new_n944), .A3(new_n886), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT105), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n903), .A2(new_n938), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n897), .B1(new_n936), .B2(new_n930), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n941), .A2(new_n952), .A3(new_n886), .A4(new_n946), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n947), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n953), .B2(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT106), .B1(new_n947), .B2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  XNOR2_X1  g539(.A(KEYINPUT107), .B(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n509), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G40), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n474), .A2(new_n481), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT109), .Z(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(G1996), .A3(new_n817), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT110), .Z(new_n973));
  NOR2_X1   g548(.A1(new_n701), .A2(new_n691), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n754), .B(G2067), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n970), .A2(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT108), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n975), .A2(new_n971), .B1(new_n977), .B2(new_n818), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n754), .A2(G2067), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n971), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n977), .B(KEYINPUT46), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n975), .A2(new_n971), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n971), .A2(new_n817), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n973), .A2(new_n978), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n701), .B(new_n691), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n971), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n970), .A2(G1986), .A3(G290), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT48), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n985), .A2(new_n990), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT114), .B(G1981), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G86), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n583), .B1(new_n526), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n517), .B1(new_n578), .B2(new_n579), .ZN(new_n1002));
  OAI21_X1  g577(.A(G1981), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1003), .A3(KEYINPUT115), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND3_X1  g580(.A1(G305), .A2(new_n1005), .A3(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n485), .A2(G126), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n460), .B1(new_n1013), .B2(new_n499), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n464), .A2(new_n485), .A3(new_n497), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n495), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT4), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n470), .A2(new_n471), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n503), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1012), .B1(new_n968), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1004), .A2(new_n1008), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1011), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT117), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1011), .A2(new_n1022), .A3(new_n1026), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G288), .A2(G1976), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1028), .A2(new_n1029), .B1(new_n723), .B2(new_n998), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1022), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n576), .A2(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1022), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1384), .ZN(new_n1036));
  INV_X1    g611(.A(new_n503), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT4), .B1(new_n629), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n499), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n485), .B2(G126), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n495), .B(new_n1015), .C1(new_n1040), .C2(new_n460), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1036), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n1043));
  INV_X1    g618(.A(new_n473), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n629), .B2(G125), .ZN(new_n1045));
  OAI211_X1 g620(.A(G40), .B(new_n1043), .C1(new_n1045), .C2(new_n464), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1033), .B(G8), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1032), .B1(new_n576), .B2(G1976), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1028), .A2(new_n1035), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n1052), .B(KEYINPUT55), .Z(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1046), .B1(new_n1021), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1042), .A2(new_n1058), .A3(KEYINPUT50), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1056), .B(new_n1057), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT45), .B(new_n965), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n509), .A2(KEYINPUT111), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1046), .B1(new_n969), .B2(new_n1042), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1971), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(G8), .B(new_n1053), .C1(new_n1062), .C2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1030), .A2(new_n1031), .B1(new_n1051), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1067), .A2(new_n1068), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n559), .A2(new_n563), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1075), .B(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(G160), .B(G40), .C1(new_n1042), .C2(KEYINPUT50), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1021), .A2(new_n1055), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n771), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1074), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1074), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(KEYINPUT61), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1091));
  INV_X1    g666(.A(G1348), .ZN(new_n1092));
  INV_X1    g667(.A(G2067), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1046), .A2(new_n1042), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(KEYINPUT60), .B2(new_n606), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n1102), .C1(new_n1046), .C2(new_n1042), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1996), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1067), .A2(new_n1108), .A3(new_n1068), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1107), .A2(KEYINPUT122), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT122), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1101), .B1(new_n1112), .B2(new_n550), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1110), .A2(new_n1111), .A3(new_n853), .A4(new_n1100), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1090), .B(new_n1099), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1095), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n606), .A3(new_n1088), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1087), .A3(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1079), .A2(new_n1080), .A3(G2090), .ZN(new_n1119));
  OAI21_X1  g694(.A(G8), .B1(new_n1069), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1053), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1070), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1051), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1067), .A2(new_n747), .A3(new_n1068), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1961), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1091), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1046), .B1(new_n966), .B2(new_n969), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(G2078), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1067), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1128), .A2(new_n1127), .B1(new_n1091), .B2(new_n1130), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1068), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(G301), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(KEYINPUT54), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1124), .A2(new_n1126), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1135), .A2(G171), .ZN(new_n1144));
  AOI21_X1  g719(.A(G301), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1068), .A2(new_n1138), .ZN(new_n1147));
  INV_X1    g722(.A(new_n796), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1056), .B(new_n828), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(G168), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(G8), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1153));
  AOI21_X1  g728(.A(G168), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1151), .B(G8), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1146), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1142), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1071), .B1(new_n1118), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1034), .B(new_n1049), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT50), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1046), .B1(new_n1021), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1164), .B(new_n1057), .C1(new_n1021), .C2(new_n1055), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n968), .B1(new_n1021), .B2(KEYINPUT45), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1167), .B2(G1971), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1053), .B1(new_n1168), .B2(G8), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1162), .B1(new_n1169), .B2(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1122), .B2(new_n1070), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(G8), .A3(G168), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1161), .B1(new_n1175), .B2(KEYINPUT63), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT119), .B(new_n1177), .C1(new_n1178), .C2(new_n1174), .ZN(new_n1179));
  OAI21_X1  g754(.A(G8), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1051), .B1(new_n1121), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1174), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(KEYINPUT63), .A3(new_n1070), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1176), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1153), .A2(new_n1156), .A3(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n1124), .A3(new_n1126), .A4(new_n1145), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT125), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1145), .A4(new_n1186), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1157), .A2(KEYINPUT62), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1160), .A2(new_n1184), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  XNOR2_X1  g770(.A(G290), .B(new_n736), .ZN(new_n1196));
  OR2_X1    g771(.A1(new_n1196), .A2(new_n970), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n993), .A2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1195), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n997), .B1(new_n1199), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g776(.A(new_n667), .B1(new_n650), .B2(new_n651), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n885), .B2(new_n886), .ZN(new_n1204));
  INV_X1    g778(.A(G229), .ZN(new_n1205));
  AND4_X1   g779(.A1(G319), .A2(new_n957), .A3(new_n1204), .A4(new_n1205), .ZN(G308));
  NAND4_X1  g780(.A1(new_n957), .A2(new_n1204), .A3(G319), .A4(new_n1205), .ZN(G225));
endmodule


