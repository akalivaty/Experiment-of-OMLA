//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT75), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n197), .C1(G119), .C2(new_n196), .ZN(new_n198));
  XNOR2_X1  g012(.A(G119), .B(G128), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  AOI22_X1  g014(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT16), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n206), .A2(G146), .A3(new_n207), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n201), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n207), .A3(G146), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(G146), .ZN(new_n213));
  XNOR2_X1  g027(.A(G125), .B(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n192), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n191), .A2(new_n210), .A3(new_n216), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G217), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G234), .B2(new_n221), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT74), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n220), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n221), .B1(new_n225), .B2(G234), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n234), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n239), .A3(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n196), .B1(new_n243), .B2(KEYINPUT69), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT1), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT66), .B1(new_n236), .B2(G143), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n237), .A2(new_n239), .A3(new_n251), .A4(G143), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT1), .B(new_n196), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n233), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n248), .B1(new_n213), .B2(G143), .ZN(new_n256));
  AND4_X1   g070(.A1(new_n251), .A2(new_n237), .A3(new_n239), .A4(G143), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n255), .B(G128), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT1), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n245), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(new_n196), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT71), .B(new_n258), .C1(new_n261), .C2(new_n241), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G137), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n265), .B2(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT11), .B1(new_n267), .B2(G134), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n267), .A2(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(KEYINPUT68), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(new_n267), .A3(KEYINPUT11), .A4(G134), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n271), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n273), .B2(new_n265), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n254), .A2(new_n262), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n194), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G119), .ZN(new_n284));
  INV_X1    g098(.A(G113), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(KEYINPUT2), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(KEYINPUT2), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n282), .B(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n284), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT2), .B(G113), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n291), .A3(KEYINPUT70), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n268), .B(new_n263), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(new_n276), .ZN(new_n298));
  OAI21_X1  g112(.A(G131), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n277), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT0), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n196), .A3(KEYINPUT64), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(KEYINPUT0), .B2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n240), .A2(new_n234), .ZN(new_n307));
  INV_X1    g121(.A(new_n235), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n196), .B1(new_n250), .B2(new_n252), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(KEYINPUT0), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n296), .B1(new_n300), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n281), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n300), .A2(new_n311), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n295), .B1(new_n281), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI211_X1 g131(.A(KEYINPUT73), .B(new_n295), .C1(new_n281), .C2(new_n314), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT28), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT28), .B1(new_n281), .B2(new_n312), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT27), .Z(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n320), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(G902), .B1(new_n319), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G128), .A3(new_n246), .ZN(new_n332));
  INV_X1    g146(.A(new_n241), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n332), .A2(new_n333), .B1(new_n255), .B2(new_n310), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n314), .B1(new_n334), .B2(new_n279), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n295), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n300), .B2(new_n311), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n281), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n337), .A2(new_n339), .B1(new_n281), .B2(new_n312), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n321), .B1(new_n340), .B2(new_n326), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n296), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n313), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(new_n320), .A3(new_n327), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n330), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n313), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n327), .ZN(new_n349));
  INV_X1    g163(.A(new_n320), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n281), .A2(new_n312), .B1(new_n335), .B2(new_n296), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n350), .B(new_n326), .C1(new_n351), .C2(new_n342), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n352), .A4(new_n321), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n329), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(G472), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT32), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n281), .A2(new_n338), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n258), .B1(new_n261), .B2(new_n241), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n358), .A2(new_n280), .B1(new_n300), .B2(new_n311), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n296), .B1(new_n359), .B2(KEYINPUT30), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n313), .B(new_n326), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n340), .A2(KEYINPUT31), .A3(new_n326), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n350), .B1(new_n351), .B2(new_n342), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n363), .A2(new_n364), .B1(new_n365), .B2(new_n327), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n356), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n327), .ZN(new_n370));
  AND4_X1   g184(.A1(KEYINPUT31), .A2(new_n347), .A3(new_n313), .A4(new_n326), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT31), .B1(new_n340), .B2(new_n326), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT32), .A3(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n232), .B1(new_n355), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT9), .B(G234), .ZN(new_n377));
  OAI21_X1  g191(.A(G221), .B1(new_n377), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT78), .B(G469), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n300), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT77), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(G107), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n384), .B2(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n389), .A2(new_n392), .A3(new_n393), .A4(new_n385), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n334), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G128), .B1(new_n235), .B2(new_n255), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n250), .A2(new_n252), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n258), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n383), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT12), .ZN(new_n402));
  INV_X1    g216(.A(new_n395), .ZN(new_n403));
  INV_X1    g217(.A(new_n399), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n253), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT10), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT76), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n400), .B2(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n395), .A2(new_n406), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n254), .A2(new_n262), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n389), .A2(new_n392), .A3(new_n385), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(G101), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n311), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n410), .A2(new_n412), .A3(new_n382), .A4(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT12), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n383), .C1(new_n397), .C2(new_n400), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G140), .ZN(new_n423));
  INV_X1    g237(.A(G227), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G953), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n402), .A2(new_n420), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT76), .B1(new_n405), .B2(new_n406), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n400), .A2(new_n408), .A3(KEYINPUT10), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n419), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n412), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n300), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n427), .B1(new_n433), .B2(new_n420), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT79), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n420), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n407), .A2(new_n409), .B1(new_n311), .B2(new_n418), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n382), .B1(new_n438), .B2(new_n412), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n435), .B(new_n426), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n221), .B(new_n381), .C1(new_n436), .C2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n437), .A2(new_n426), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n402), .A2(new_n420), .A3(new_n422), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n443), .A2(new_n433), .B1(new_n444), .B2(new_n426), .ZN(new_n445));
  OAI21_X1  g259(.A(G469), .B1(new_n445), .B2(G902), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n379), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n187), .A2(G224), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT80), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT81), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n247), .A2(G125), .A3(new_n253), .ZN(new_n456));
  INV_X1    g270(.A(new_n309), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT0), .B(G128), .C1(new_n256), .C2(new_n257), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n204), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n455), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n204), .B(new_n258), .C1(new_n261), .C2(new_n241), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n463), .A3(new_n454), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n415), .A2(new_n292), .A3(new_n294), .A4(new_n417), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G122), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT5), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(G113), .C1(KEYINPUT5), .C2(new_n282), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n403), .A2(new_n288), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT6), .ZN(new_n473));
  INV_X1    g287(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n474), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n465), .A2(new_n466), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n453), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n461), .B2(new_n463), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n468), .B(new_n483), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n288), .A2(new_n470), .A3(new_n394), .A4(new_n388), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n470), .A2(new_n288), .B1(new_n394), .B2(new_n388), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n472), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n459), .B1(new_n334), .B2(new_n204), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n490), .B2(new_n481), .ZN(new_n491));
  AND4_X1   g305(.A1(KEYINPUT84), .A2(new_n461), .A3(new_n463), .A4(new_n481), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n221), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n473), .B(new_n477), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n466), .B1(new_n495), .B2(new_n465), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n451), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n465), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n476), .A2(new_n478), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT82), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n490), .A2(KEYINPUT84), .A3(new_n481), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n461), .A2(new_n463), .A3(new_n481), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n505), .B2(new_n489), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n500), .A2(new_n506), .A3(new_n450), .A4(new_n479), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n449), .B1(new_n497), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n215), .B1(new_n236), .B2(new_n214), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n187), .A3(G214), .ZN(new_n514));
  NAND2_X1  g328(.A1(KEYINPUT85), .A2(G143), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(KEYINPUT85), .A2(G143), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(KEYINPUT85), .A2(G143), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(G214), .A3(new_n322), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n520), .C1(new_n521), .C2(new_n271), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n519), .A2(new_n515), .B1(new_n322), .B2(G214), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n514), .A2(new_n517), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n512), .B(new_n522), .C1(new_n525), .C2(new_n521), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n518), .A2(new_n271), .A3(new_n520), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n271), .B1(new_n518), .B2(new_n520), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n212), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT19), .B1(new_n214), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n214), .A2(new_n530), .A3(KEYINPUT19), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n240), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n526), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n384), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT17), .ZN(new_n540));
  INV_X1    g354(.A(new_n208), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT17), .B(G131), .C1(new_n523), .C2(new_n524), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n212), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n537), .B(new_n526), .C1(new_n540), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n511), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT20), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g361(.A(KEYINPUT87), .B(new_n511), .C1(new_n539), .C2(new_n544), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n544), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n518), .A2(new_n271), .A3(new_n520), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n525), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n533), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n531), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n212), .C1(new_n554), .C2(new_n240), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n537), .B1(new_n555), .B2(new_n526), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n510), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(KEYINPUT87), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n209), .A2(new_n208), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n560), .B(new_n542), .C1(new_n552), .C2(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n537), .B1(new_n561), .B2(new_n526), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n221), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G475), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n509), .B1(new_n549), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n539), .A2(new_n544), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n546), .B1(new_n567), .B2(new_n510), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n558), .B1(G475), .B2(new_n563), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n557), .A2(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n545), .A2(new_n546), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(KEYINPUT20), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT88), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G122), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT89), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G122), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n283), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n575), .A2(G116), .ZN(new_n580));
  OAI21_X1  g394(.A(G107), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT89), .B(G122), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n391), .B(new_n582), .C1(new_n583), .C2(new_n283), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n234), .A2(G128), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n196), .A2(G143), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n264), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n196), .B2(G143), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n234), .A2(KEYINPUT13), .A3(G128), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n587), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n592), .A2(new_n593), .A3(G134), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n592), .B2(G134), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n585), .B(new_n588), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT14), .B1(new_n583), .B2(new_n283), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(G107), .C1(new_n580), .C2(new_n579), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n264), .B1(new_n586), .B2(new_n587), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(KEYINPUT91), .A3(new_n588), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n602));
  INV_X1    g416(.A(new_n588), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n599), .ZN(new_n604));
  OAI221_X1 g418(.A(new_n582), .B1(KEYINPUT14), .B2(new_n391), .C1(new_n583), .C2(new_n283), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n598), .A2(new_n601), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n377), .A2(new_n225), .A3(G953), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n606), .A3(new_n608), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n221), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n613), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n574), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n187), .A2(G952), .ZN(new_n619));
  NAND2_X1  g433(.A1(G234), .A2(G237), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(G902), .A3(G953), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT92), .Z(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n447), .A2(new_n508), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n376), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n393), .ZN(G3));
  OR2_X1    g445(.A1(new_n228), .A2(new_n231), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n373), .B2(new_n221), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n366), .A2(new_n368), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n447), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT93), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n596), .A2(new_n606), .A3(new_n639), .A4(new_n608), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n610), .A2(KEYINPUT33), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT94), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n612), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n607), .B2(new_n609), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n642), .A3(new_n648), .A4(new_n640), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n614), .A2(G902), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n644), .A2(new_n646), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n613), .A2(new_n614), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n574), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n508), .A3(new_n626), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT95), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n655), .A2(new_n508), .A3(new_n658), .A4(new_n626), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n638), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NOR2_X1   g477(.A1(new_n549), .A2(new_n565), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n626), .A3(new_n616), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT96), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n497), .A2(new_n507), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n448), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n638), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT97), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n634), .A2(new_n635), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(new_n217), .Z(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n230), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n224), .B2(new_n227), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n675), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT99), .A4(new_n680), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n629), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT37), .B(G110), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  OAI21_X1  g500(.A(new_n621), .B1(G900), .B2(new_n624), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n616), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n508), .A2(new_n681), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n690), .B(new_n447), .C1(new_n355), .C2(new_n375), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n366), .A2(new_n356), .A3(new_n368), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT32), .B1(new_n373), .B2(new_n367), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n354), .A2(G472), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(KEYINPUT100), .A3(new_n447), .A4(new_n690), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XNOR2_X1  g515(.A(new_n687), .B(KEYINPUT39), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n447), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n348), .A2(new_n326), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n221), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n317), .A2(new_n326), .A3(new_n318), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n369), .A2(new_n374), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n574), .A2(new_n617), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n667), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n448), .A3(new_n680), .ZN(new_n715));
  OR4_X1    g529(.A1(new_n704), .A2(new_n705), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n566), .A2(new_n653), .A3(new_n573), .A4(new_n687), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n668), .B2(new_n720), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n566), .A2(new_n653), .A3(new_n573), .A4(new_n687), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n508), .A3(KEYINPUT102), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n447), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n681), .B1(new_n355), .B2(new_n375), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n718), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n680), .B1(new_n696), .B2(new_n697), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n722), .A2(new_n508), .A3(KEYINPUT102), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT102), .B1(new_n722), .B2(new_n508), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n730), .A3(KEYINPUT103), .A4(new_n447), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(G469), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n426), .B1(new_n437), .B2(new_n439), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT79), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n440), .A3(new_n428), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n734), .B(new_n735), .C1(new_n738), .C2(new_n221), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n221), .B1(new_n436), .B2(new_n441), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT104), .B1(new_n740), .B2(G469), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n378), .B(new_n442), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n632), .B1(new_n696), .B2(new_n697), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n660), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n669), .A3(new_n744), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NOR2_X1   g563(.A1(new_n742), .A2(new_n668), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n628), .A3(new_n727), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  XNOR2_X1  g566(.A(KEYINPUT105), .B(G472), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n366), .B2(G902), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n326), .B1(new_n319), .B2(new_n350), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n371), .A2(new_n372), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n367), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n757), .A3(new_n232), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n711), .A2(new_n508), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n627), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n743), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT106), .B(G122), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G24));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n757), .A3(new_n681), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT107), .A4(new_n681), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n720), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n750), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NAND2_X1  g584(.A1(new_n442), .A2(new_n446), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n667), .A2(new_n449), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n378), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n447), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n774), .A2(new_n744), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n720), .A2(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n695), .B1(G472), .B2(new_n354), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n374), .A2(KEYINPUT109), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n694), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n232), .A3(new_n722), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n774), .A2(new_n776), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n271), .ZN(G33));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n689), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OR2_X1    g605(.A1(new_n445), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n445), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT110), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n798), .B(new_n442), .C1(new_n797), .C2(new_n796), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT110), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n379), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n702), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT43), .B1(new_n574), .B2(new_n653), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n574), .B(KEYINPUT112), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n654), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n808), .B2(KEYINPUT43), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n809), .A2(new_n676), .A3(new_n680), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT44), .Z(new_n811));
  XOR2_X1   g625(.A(new_n772), .B(KEYINPUT113), .Z(new_n812));
  NAND3_X1  g626(.A1(new_n805), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G137), .ZN(G39));
  XOR2_X1   g628(.A(new_n802), .B(KEYINPUT47), .Z(new_n815));
  NAND3_X1  g629(.A1(new_n772), .A2(new_n632), .A3(new_n722), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n698), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND4_X1  g633(.A1(new_n808), .A2(new_n232), .A3(new_n378), .A4(new_n448), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n710), .A3(new_n714), .ZN(new_n821));
  INV_X1    g635(.A(new_n442), .ZN(new_n822));
  INV_X1    g636(.A(new_n741), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n740), .A2(KEYINPUT104), .A3(G469), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n821), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n617), .A2(new_n664), .A3(new_n687), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n725), .A2(new_n773), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n786), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n768), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n654), .A2(new_n566), .A3(new_n573), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n508), .A2(new_n618), .A3(new_n626), .A4(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n637), .A2(new_n836), .B1(new_n376), .B2(new_n629), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n684), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n838), .A3(new_n790), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n751), .A2(new_n748), .A3(new_n745), .A4(new_n761), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(new_n788), .A3(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n726), .A2(new_n731), .B1(new_n693), .B2(new_n699), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n710), .A2(new_n680), .A3(new_n687), .A4(new_n711), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n447), .A2(new_n508), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n750), .B2(new_n768), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n732), .A3(new_n700), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n830), .A2(new_n841), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n843), .A2(new_n847), .A3(new_n700), .A4(new_n732), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n843), .B1(new_n842), .B2(new_n847), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n850), .A2(KEYINPUT114), .A3(new_n848), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n841), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n851), .B1(KEYINPUT53), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n830), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n850), .A2(new_n848), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n823), .A2(new_n824), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n378), .A3(new_n442), .A4(new_n508), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n727), .A2(new_n628), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n748), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n745), .A2(new_n761), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n783), .A2(new_n781), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n632), .B1(new_n868), .B2(new_n780), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n722), .A3(new_n774), .A4(new_n776), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n870), .A2(KEYINPUT42), .B1(new_n777), .B2(new_n778), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(KEYINPUT53), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n839), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n860), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n859), .B(KEYINPUT115), .C1(KEYINPUT54), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(KEYINPUT115), .B2(new_n859), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n809), .A2(new_n621), .ZN(new_n880));
  INV_X1    g694(.A(new_n758), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n882), .A2(new_n448), .A3(new_n714), .A4(new_n742), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT50), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n742), .A2(new_n449), .A3(new_n667), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n710), .A2(new_n632), .A3(new_n621), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n574), .A3(new_n654), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n766), .A2(new_n767), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n885), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n884), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n882), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n812), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n825), .A2(new_n379), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n815), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n897));
  INV_X1    g711(.A(new_n869), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT48), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n885), .A2(new_n655), .A3(new_n886), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n619), .B(new_n901), .C1(new_n882), .C2(new_n863), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n879), .A2(new_n896), .A3(new_n897), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n829), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n187), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n857), .A2(new_n830), .B1(new_n873), .B2(new_n875), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n221), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n499), .B(KEYINPUT117), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n465), .B(KEYINPUT55), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n912), .B(new_n913), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n909), .B2(new_n221), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n451), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(G51));
  OR2_X1    g739(.A1(new_n920), .A2(new_n794), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(KEYINPUT120), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n877), .B(KEYINPUT54), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n795), .B(KEYINPUT57), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n926), .A2(KEYINPUT120), .B1(new_n738), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n907), .B1(new_n927), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n544), .A3(new_n539), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .A4(new_n567), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n908), .A3(new_n935), .ZN(G60));
  NAND3_X1  g750(.A1(new_n644), .A2(new_n646), .A3(new_n649), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n879), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n907), .B1(new_n928), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(G63));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n877), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n909), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n952), .A3(new_n229), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n950), .A2(new_n952), .A3(new_n955), .A4(new_n229), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n678), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT122), .B1(new_n877), .B2(new_n949), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n909), .A2(new_n951), .A3(new_n948), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(KEYINPUT61), .A3(new_n908), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n946), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n678), .B1(new_n950), .B2(new_n952), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n907), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n954), .A4(new_n956), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n961), .A2(new_n908), .A3(new_n953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n965), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n622), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n867), .A2(new_n838), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n975), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n912), .B1(G898), .B2(new_n187), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  OAI21_X1  g792(.A(new_n339), .B1(KEYINPUT30), .B2(new_n359), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n554), .ZN(new_n980));
  INV_X1    g794(.A(G900), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n187), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n842), .A2(new_n769), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n871), .A2(new_n984), .A3(new_n790), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n818), .A2(new_n813), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n898), .A2(new_n759), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n805), .A2(KEYINPUT126), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n805), .A2(new_n988), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n987), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n982), .B1(new_n993), .B2(new_n187), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n818), .A2(new_n813), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n984), .A2(new_n716), .A3(new_n985), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n772), .A2(new_n618), .A3(new_n835), .ZN(new_n999));
  OR3_X1    g813(.A1(new_n376), .A2(new_n703), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n995), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n980), .B1(new_n1001), .B2(new_n187), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n994), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n349), .B2(new_n361), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n907), .B1(new_n858), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1009), .B1(new_n993), .B2(new_n975), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n340), .A2(new_n327), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1008), .B1(new_n1001), .B2(new_n974), .ZN(new_n1015));
  INV_X1    g829(.A(new_n706), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1015), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1014), .B1(new_n1018), .B2(new_n1020), .ZN(G57));
endmodule


