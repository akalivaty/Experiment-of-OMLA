//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G221), .A2(G219), .A3(G218), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT69), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT71), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g051(.A(G137), .B(new_n466), .C1(new_n469), .C2(new_n470), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n466), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(new_n466), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n464), .A2(new_n466), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AOI211_X1 g066(.A(new_n485), .B(new_n488), .C1(new_n491), .C2(G136), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n466), .B2(G114), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n469), .B2(new_n470), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n464), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n466), .C1(new_n469), .C2(new_n470), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n464), .A2(new_n507), .A3(G138), .A4(new_n466), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(G75), .B2(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(KEYINPUT75), .A3(G62), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n512), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n513), .A2(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G88), .B1(new_n526), .B2(G50), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n520), .A2(new_n528), .ZN(G166));
  AOI22_X1  g104(.A1(new_n524), .A2(G89), .B1(new_n526), .B2(G51), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n536), .A2(new_n532), .A3(new_n534), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  XOR2_X1   g118(.A(KEYINPUT77), .B(G52), .Z(new_n544));
  AOI22_X1  g119(.A1(new_n524), .A2(G90), .B1(new_n526), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT5), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G64), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n512), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n545), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n515), .A2(G56), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n512), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  NOR2_X1   g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n547), .A2(new_n546), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(G543), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n546), .A2(new_n547), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n557), .A2(new_n558), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n576), .A2(G53), .A3(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(new_n523), .ZN(new_n579));
  INV_X1    g154(.A(new_n577), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  OAI211_X1 g159(.A(G53), .B(G543), .C1(new_n557), .C2(new_n558), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT9), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n583), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n574), .B1(new_n587), .B2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G166), .ZN(G303));
  NAND2_X1  g165(.A1(new_n524), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(G49), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n571), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n524), .A2(G86), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n512), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n559), .A2(new_n604), .B1(new_n561), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n561), .B2(KEYINPUT81), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n526), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(G66), .B1(new_n546), .B2(new_n547), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n613), .A2(new_n615), .B1(new_n618), .B2(G651), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n559), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n515), .A2(new_n579), .A3(KEYINPUT10), .A4(G92), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n611), .B1(new_n625), .B2(G868), .ZN(G284));
  XOR2_X1   g201(.A(G284), .B(KEYINPUT82), .Z(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(new_n574), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n575), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n586), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT79), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n578), .A2(new_n582), .B1(KEYINPUT9), .B2(new_n585), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n584), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n629), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n628), .B1(new_n636), .B2(G868), .ZN(G297));
  OAI21_X1  g212(.A(new_n628), .B1(new_n636), .B2(G868), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n625), .B1(new_n639), .B2(G860), .ZN(G148));
  NOR2_X1   g215(.A1(new_n564), .A2(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n625), .A2(new_n639), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n486), .A2(G123), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n491), .A2(G135), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2096), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(G2096), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n464), .A2(new_n478), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT13), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2451), .B(G2454), .Z(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(G14), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT87), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT17), .Z(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT90), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n682), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n686));
  INV_X1    g261(.A(new_n678), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n680), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n680), .A2(new_n681), .A3(new_n678), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT18), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n684), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n706), .B(new_n705), .S(new_n698), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G229));
  NAND2_X1  g290(.A1(new_n491), .A2(G131), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G107), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(new_n721), .B1(G119), .B2(new_n486), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n716), .A2(KEYINPUT92), .A3(new_n722), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n725), .A2(G29), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G25), .B2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(G290), .A2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G24), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT93), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1986), .Z(new_n737));
  AND3_X1   g312(.A1(new_n730), .A2(new_n731), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(G6), .ZN(new_n739));
  INV_X1    g314(.A(G305), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT94), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT32), .B(G1981), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n733), .A2(G23), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n594), .B2(new_n733), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT33), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1976), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G22), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G166), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1971), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n742), .A2(new_n744), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n745), .A2(new_n749), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n755));
  OAI21_X1  g330(.A(new_n738), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT36), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n754), .A2(new_n755), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n755), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n738), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n733), .A2(G5), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G301), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n564), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G16), .B2(G19), .ZN(new_n769));
  INV_X1    g344(.A(G1341), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G29), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n651), .A2(new_n772), .B1(new_n766), .B2(new_n765), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n733), .A2(G21), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G168), .B2(new_n733), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n771), .B(new_n773), .C1(new_n776), .C2(G1966), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(KEYINPUT24), .B2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(KEYINPUT24), .B2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n481), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2084), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n772), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n491), .A2(G140), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  INV_X1    g362(.A(G116), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G2105), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n486), .B2(G128), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(G29), .ZN(new_n792));
  AOI211_X1 g367(.A(KEYINPUT96), .B(new_n772), .C1(new_n786), .C2(new_n790), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n784), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n625), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G4), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n776), .B2(G1966), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n782), .A2(new_n795), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n733), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n636), .B2(new_n733), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT100), .B(G1956), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n772), .A2(G32), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n491), .A2(G141), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n478), .A2(G105), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT26), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n811), .B(new_n813), .C1(G129), .C2(new_n486), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n809), .B1(new_n816), .B2(new_n772), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT27), .B(G1996), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  NAND2_X1  g396(.A1(G162), .A2(G29), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G29), .B2(G35), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT29), .B(G2090), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT25), .Z(new_n828));
  AOI22_X1  g403(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n466), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n491), .B2(G139), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G29), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G29), .B2(G33), .ZN(new_n833));
  INV_X1    g408(.A(G2072), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(G164), .A2(G29), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G27), .B2(G29), .ZN(new_n838));
  INV_X1    g413(.A(G2078), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n826), .A2(new_n835), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n823), .A2(new_n825), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT31), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(G11), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(G11), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT30), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(G28), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n772), .B1(new_n847), .B2(G28), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n845), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n769), .B2(new_n770), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n817), .A2(new_n819), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n842), .A2(new_n843), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n821), .A2(new_n841), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n802), .A2(new_n808), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n763), .A2(KEYINPUT102), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT102), .B1(new_n763), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(G311));
  NAND2_X1  g433(.A1(new_n763), .A2(new_n855), .ZN(G150));
  NAND2_X1  g434(.A1(new_n625), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n524), .A2(G81), .B1(new_n526), .B2(G43), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n524), .A2(G93), .B1(new_n526), .B2(G55), .ZN(new_n863));
  INV_X1    g438(.A(G56), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n513), .B2(new_n514), .ZN(new_n865));
  INV_X1    g440(.A(new_n555), .ZN(new_n866));
  OAI21_X1  g441(.A(G651), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G67), .B1(new_n546), .B2(new_n547), .ZN(new_n868));
  NAND2_X1  g443(.A1(G80), .A2(G543), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G651), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n862), .A2(new_n863), .A3(new_n867), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(G55), .B(G543), .C1(new_n557), .C2(new_n558), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n559), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n512), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n556), .A2(new_n563), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n861), .B(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(G860), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n863), .A2(new_n871), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G860), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT103), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  OR2_X1    g462(.A1(new_n883), .A2(new_n887), .ZN(G145));
  XNOR2_X1  g463(.A(G160), .B(new_n651), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G162), .ZN(new_n890));
  INV_X1    g465(.A(new_n791), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n816), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n815), .A2(new_n791), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G164), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n510), .A3(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n831), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n831), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n656), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n725), .A2(new_n726), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n491), .A2(G142), .ZN(new_n905));
  OAI21_X1  g480(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n906));
  INV_X1    g481(.A(G118), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(G2105), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n486), .B2(G130), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n904), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n656), .A3(new_n912), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n917), .A3(KEYINPUT104), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT104), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n902), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n918), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n922), .A2(new_n919), .A3(new_n901), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n890), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n917), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n890), .B1(new_n902), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n901), .B1(new_n922), .B2(new_n919), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n924), .A2(KEYINPUT40), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT40), .B1(new_n924), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(G395));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(G868), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n884), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n642), .B(new_n878), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n619), .A2(new_n624), .ZN(new_n936));
  NOR2_X1   g511(.A1(G299), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n633), .A2(new_n635), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n625), .B1(new_n938), .B2(new_n574), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n937), .B2(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(G299), .A2(new_n936), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n636), .A2(new_n625), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(new_n935), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n943), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G166), .A2(G288), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n594), .B1(new_n520), .B2(new_n528), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(new_n740), .ZN(new_n958));
  OAI211_X1 g533(.A(G305), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n955), .A2(new_n958), .A3(new_n956), .A4(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n954), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G868), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n952), .B2(new_n954), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n934), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(new_n932), .A3(G868), .A4(new_n965), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(G295));
  AND2_X1   g546(.A1(new_n968), .A2(new_n970), .ZN(G331));
  NAND4_X1  g547(.A1(new_n530), .A2(new_n545), .A3(new_n541), .A4(new_n551), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n515), .A2(new_n540), .ZN(new_n974));
  INV_X1    g549(.A(new_n539), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n536), .B1(new_n532), .B2(new_n534), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G89), .ZN(new_n978));
  INV_X1    g553(.A(G51), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n559), .A2(new_n978), .B1(new_n561), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G90), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT77), .B(G52), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n559), .A2(new_n981), .B1(new_n561), .B2(new_n982), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n977), .A2(new_n980), .B1(new_n983), .B2(new_n550), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n878), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n973), .A2(new_n872), .A3(new_n984), .A4(new_n877), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n945), .A2(new_n948), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(KEYINPUT108), .A3(new_n987), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n879), .A2(new_n991), .A3(new_n984), .A4(new_n973), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n940), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n963), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(new_n994), .A3(new_n963), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n997), .ZN(new_n1002));
  INV_X1    g577(.A(new_n963), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n945), .A2(new_n948), .A3(new_n992), .A4(new_n990), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n940), .A2(new_n987), .A3(new_n986), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1000), .B(KEYINPUT44), .C1(new_n1001), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n995), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1003), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(new_n1001), .A3(new_n997), .A4(new_n998), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT110), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT109), .B1(new_n999), .B2(KEYINPUT43), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT110), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1008), .B1(new_n1018), .B2(new_n1022), .ZN(G397));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n510), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n477), .A2(new_n479), .A3(G40), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n467), .A2(new_n475), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n729), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n904), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2067), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n791), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1996), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n815), .B(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(G290), .B(G1986), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1030), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1026), .A2(G1384), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1029), .B1(new_n510), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1027), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1045), .B2(G2078), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n467), .A2(new_n475), .A3(new_n1028), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n510), .A2(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n504), .B2(new_n509), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(KEYINPUT45), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n1053));
  NOR2_X1   g628(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n510), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1047), .B(new_n1055), .C1(new_n1056), .C2(new_n1050), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n766), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1046), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n473), .A2(KEYINPUT121), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n466), .B1(new_n473), .B2(KEYINPUT121), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1027), .A2(new_n1064), .A3(new_n1048), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1046), .A2(G301), .A3(new_n1058), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1041), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(new_n1072), .C1(new_n1071), .C2(G288), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT112), .B(G86), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n599), .B1(new_n559), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1076), .A2(G1981), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G305), .A2(G1981), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(G1981), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1070), .A3(new_n1081), .ZN(new_n1082));
  OAI221_X1 g657(.A(G8), .B1(new_n1071), .B2(G288), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT52), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1057), .A2(G2090), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1971), .B1(new_n1044), .B2(new_n1027), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT55), .B(G8), .C1(new_n520), .C2(new_n528), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G166), .B2(new_n1069), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(G8), .C1(new_n1088), .C2(new_n1087), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1086), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1067), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1966), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1103));
  INV_X1    g678(.A(G2084), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1047), .A4(new_n1055), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(G168), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  AND2_X1   g682(.A1(KEYINPUT118), .A2(G8), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(G286), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1107), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT119), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1111), .A4(new_n1109), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1046), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(KEYINPUT54), .C1(G171), .C2(new_n1059), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1100), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1052), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1057), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1057), .B2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n636), .A2(KEYINPUT57), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n629), .B2(new_n634), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1057), .A2(new_n1126), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT113), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1057), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1138), .A2(new_n1139), .B1(new_n1052), .B2(new_n1123), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1140), .B2(new_n1133), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1133), .B(new_n1124), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(KEYINPUT115), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1135), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1068), .A2(new_n1033), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1057), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT60), .B(new_n1147), .C1(new_n1148), .C2(G1348), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1149), .A2(KEYINPUT117), .A3(new_n936), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n936), .B1(new_n1149), .B2(KEYINPUT117), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1150), .A2(new_n1151), .B1(KEYINPUT117), .B2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1148), .B2(G1348), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(KEYINPUT60), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1135), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1129), .A2(KEYINPUT116), .A3(new_n1134), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(KEYINPUT61), .A3(new_n1158), .A4(new_n1142), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT58), .B(G1341), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1045), .A2(G1996), .B1(new_n1068), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n564), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT59), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1146), .A2(new_n1155), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1153), .A2(new_n625), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1157), .A2(new_n1165), .A3(new_n1158), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1122), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1114), .A2(new_n1117), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1099), .A2(new_n1060), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G288), .A2(G1976), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1078), .B1(new_n1082), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1070), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1098), .A2(new_n1085), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1069), .B(G286), .C1(new_n1102), .C2(new_n1105), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1086), .A2(new_n1096), .A3(new_n1098), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1177), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1173), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1040), .B1(new_n1168), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1037), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1187), .B2(new_n1037), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(G2067), .B2(new_n791), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1030), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1030), .A2(KEYINPUT46), .A3(new_n1035), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT123), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT46), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1034), .A2(new_n816), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1030), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1198));
  AOI21_X1  g773(.A(KEYINPUT124), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1199));
  NOR2_X1   g774(.A1(G290), .A2(G1986), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1030), .A2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT126), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1201), .B(new_n1203), .Z(new_n1204));
  NOR2_X1   g779(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1038), .A2(KEYINPUT124), .A3(new_n1030), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1191), .A2(new_n1198), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT127), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1185), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g785(.A1(G227), .A2(new_n462), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n714), .A2(new_n676), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1214));
  AOI211_X1 g788(.A(new_n1213), .B(new_n1214), .C1(new_n924), .C2(new_n928), .ZN(G308));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n924), .B2(new_n928), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(new_n1016), .ZN(G225));
endmodule


