//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT69), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(new_n467), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n469), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n466), .A2(new_n477), .A3(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n462), .A2(G2104), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  INV_X1    g055(.A(G101), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G160));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT71), .Z(new_n485));
  NOR2_X1   g060(.A1(new_n472), .A2(new_n467), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n466), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n487), .A2(G124), .B1(new_n488), .B2(G136), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n485), .A2(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n470), .A2(new_n473), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n463), .A2(new_n465), .A3(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n496), .B2(new_n486), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT72), .B(KEYINPUT4), .C1(new_n496), .C2(new_n486), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT73), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT73), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT6), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n503), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n509), .B2(new_n514), .ZN(new_n518));
  AOI22_X1  g093(.A1(G50), .A2(new_n515), .B1(new_n518), .B2(G88), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n520), .B2(KEYINPUT75), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n507), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT76), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n518), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n515), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n512), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n515), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n517), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n518), .A2(G91), .B1(G651), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n505), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n559));
  NOR4_X1   g134(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT74), .A4(new_n508), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n515), .A2(KEYINPUT77), .A3(G53), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n515), .A2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n518), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  AOI22_X1  g152(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n512), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(G48), .A2(new_n515), .B1(new_n518), .B2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n518), .A2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n515), .A2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n512), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G301), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n515), .A2(G54), .B1(G651), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT80), .Z(new_n599));
  AOI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(new_n589), .ZN(G284));
  AOI21_X1  g175(.A(new_n590), .B1(new_n599), .B2(new_n589), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NOR2_X1   g182(.A1(new_n549), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n606), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(new_n495), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n480), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(G2100), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  OAI221_X1 g195(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n487), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n488), .A2(G135), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n630), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT17), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n645), .B2(new_n642), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n647), .B2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(new_n642), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n648), .A3(new_n644), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n643), .A2(new_n648), .A3(new_n645), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n665), .A3(new_n663), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n670), .C1(new_n665), .C2(new_n669), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  AND2_X1   g252(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(new_n573), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT33), .B(G1976), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n679), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(new_n687), .ZN(new_n690));
  MUX2_X1   g265(.A(G6), .B(G305), .S(G16), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT32), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n690), .A2(new_n693), .A3(KEYINPUT34), .ZN(new_n694));
  OAI221_X1 g269(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n487), .A2(G119), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n488), .A2(G131), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT85), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(G16), .A2(G24), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G290), .B2(new_n679), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n694), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n690), .A2(new_n693), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g289(.A(KEYINPUT87), .B(KEYINPUT34), .C1(new_n690), .C2(new_n693), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n678), .B(new_n709), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT25), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n466), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n721), .B(new_n723), .C1(G139), .C2(new_n488), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n728));
  INV_X1    g303(.A(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(G160), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(G32), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n487), .A2(G129), .B1(new_n488), .B2(G141), .ZN(new_n736));
  INV_X1    g311(.A(G105), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n480), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  NOR2_X1   g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(new_n732), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n725), .B2(G2072), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n727), .A2(new_n734), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n679), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n549), .B2(new_n679), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1341), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n732), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n732), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT29), .B(G2090), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n732), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  OAI221_X1 g332(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n487), .A2(G128), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G140), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n757), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n624), .A2(new_n732), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT93), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT93), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(KEYINPUT30), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n743), .B2(new_n744), .ZN(new_n774));
  AND4_X1   g349(.A1(new_n751), .A2(new_n755), .A3(new_n763), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n679), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n733), .A2(G2084), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  NOR2_X1   g358(.A1(G5), .A2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G301), .B2(new_n679), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n782), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n679), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n679), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n781), .B(new_n787), .C1(new_n789), .C2(G1966), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(G1966), .ZN(new_n791));
  NOR2_X1   g366(.A1(G164), .A2(new_n732), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G27), .B2(new_n732), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n786), .A2(new_n783), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n775), .A2(new_n779), .A3(new_n790), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n679), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n599), .B2(new_n679), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1348), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n748), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n694), .B(new_n708), .C1(new_n713), .C2(new_n715), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n717), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G67), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n517), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n515), .A2(G55), .B1(new_n507), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT97), .B(G93), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n518), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n599), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n548), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n814), .A2(new_n548), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n818), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT98), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n825), .B2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n724), .B(new_n742), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n698), .B(KEYINPUT99), .Z(new_n830));
  AOI22_X1  g405(.A1(new_n487), .A2(G130), .B1(new_n488), .B2(G142), .ZN(new_n831));
  OAI221_X1 g406(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n498), .A2(new_n499), .ZN(new_n836));
  INV_X1    g411(.A(new_n496), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT4), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n838), .A3(new_n473), .A4(new_n470), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n501), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n494), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n761), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n616), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n835), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G162), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n624), .ZN(new_n848));
  AOI21_X1  g423(.A(G37), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n846), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(new_n814), .A2(new_n589), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n609), .B(new_n822), .ZN(new_n853));
  INV_X1    g428(.A(new_n598), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n603), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n598), .A2(G299), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT41), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n857), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n853), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n573), .B(KEYINPUT101), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G290), .ZN(new_n866));
  AND2_X1   g441(.A1(G305), .A2(G303), .ZN(new_n867));
  NOR2_X1   g442(.A1(G305), .A2(G303), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT102), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT102), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n864), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n852), .B1(new_n875), .B2(new_n589), .ZN(G295));
  OAI21_X1  g451(.A(new_n852), .B1(new_n875), .B2(new_n589), .ZN(G331));
  INV_X1    g452(.A(new_n821), .ZN(new_n878));
  AOI21_X1  g453(.A(G301), .B1(new_n878), .B2(new_n819), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n820), .A2(new_n821), .A3(G171), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n882), .A3(G168), .ZN(new_n883));
  OAI21_X1  g458(.A(G286), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n883), .B(new_n884), .C1(new_n858), .C2(new_n860), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n879), .A2(new_n881), .A3(G286), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n863), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n873), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n873), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n888), .A2(KEYINPUT103), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n857), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n859), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n855), .A2(new_n856), .A3(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n898), .A2(new_n883), .A3(new_n884), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n857), .B1(new_n883), .B2(new_n884), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n873), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n891), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n895), .B1(KEYINPUT43), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n890), .A2(new_n888), .A3(new_n885), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n910), .A2(new_n893), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n891), .A2(new_n915), .A3(new_n911), .A4(new_n893), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n908), .B1(new_n906), .B2(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n909), .B1(new_n920), .B2(new_n921), .ZN(G397));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(G1384), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n842), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(KEYINPUT107), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(KEYINPUT107), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT45), .ZN(new_n928));
  INV_X1    g503(.A(G40), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n476), .A2(new_n482), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT108), .ZN(new_n932));
  INV_X1    g507(.A(G2067), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n761), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n742), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n701), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n698), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n931), .A2(G1996), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n742), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n931), .ZN(new_n945));
  XNOR2_X1  g520(.A(G290), .B(G1986), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1966), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n842), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n840), .B2(new_n841), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n930), .B1(new_n953), .B2(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n948), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G160), .A2(G40), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G2084), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT119), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n955), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(G168), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n962), .A2(G8), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  INV_X1    g550(.A(new_n965), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n964), .B1(new_n955), .B2(new_n961), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G286), .A2(G8), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n966), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n978), .A2(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT120), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n956), .B1(new_n950), .B2(new_n951), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n989), .B2(G2078), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n958), .A2(new_n960), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n783), .ZN(new_n992));
  INV_X1    g567(.A(new_n476), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT124), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n482), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n929), .B(new_n996), .C1(new_n482), .C2(new_n994), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n988), .A2(new_n993), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n990), .B(new_n992), .C1(new_n928), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G171), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n952), .A2(new_n954), .A3(new_n996), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n992), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1001), .B2(new_n992), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n990), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT54), .B(new_n1000), .C1(new_n1005), .C2(G171), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n989), .A2(new_n688), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT111), .B(G2090), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n958), .A2(new_n960), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n968), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n930), .B1(new_n953), .B2(new_n957), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  NOR2_X1   g591(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n842), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1017), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT112), .B(new_n1019), .C1(new_n840), .C2(new_n841), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1008), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1007), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n1023), .B2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n950), .A2(new_n956), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n968), .ZN(new_n1031));
  OR2_X1    g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n681), .A2(G1976), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n574), .A2(new_n1038), .A3(new_n575), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1031), .A2(new_n1039), .A3(new_n1040), .A4(new_n1035), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1034), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1014), .A2(new_n1024), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1006), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n999), .A2(G171), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(G171), .B2(new_n1005), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n985), .B(new_n1044), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT61), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n987), .A2(new_n988), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1021), .B2(G1956), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n565), .A2(new_n1053), .A3(new_n568), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n565), .B2(new_n568), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1956), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT112), .B1(G164), .B2(new_n1019), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n842), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(new_n1015), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(new_n1056), .A3(new_n1051), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT116), .ZN(new_n1065));
  INV_X1    g640(.A(new_n957), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(G164), .B2(G1384), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(new_n1060), .A3(new_n930), .A4(new_n1061), .ZN(new_n1068));
  AOI211_X1 g643(.A(new_n951), .B(new_n923), .C1(new_n840), .C2(new_n841), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n954), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1059), .A2(new_n1068), .B1(new_n1070), .B2(new_n1050), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1056), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1058), .A2(new_n1065), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1058), .A2(new_n1065), .A3(new_n1073), .A4(KEYINPUT117), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1071), .B2(new_n1056), .ZN(new_n1081));
  AND4_X1   g656(.A1(new_n1080), .A2(new_n1063), .A3(new_n1056), .A4(new_n1051), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n950), .A2(new_n951), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(new_n935), .A3(new_n930), .A4(new_n988), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n987), .A2(new_n1087), .A3(new_n935), .A4(new_n988), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n950), .B2(new_n956), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n549), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT115), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1091), .B(new_n549), .C1(KEYINPUT115), .C2(new_n1093), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1083), .A2(new_n1049), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1078), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1078), .A2(new_n1097), .A3(KEYINPUT118), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n991), .A2(new_n1102), .B1(new_n933), .B2(new_n1030), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(new_n854), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(KEYINPUT60), .B2(new_n1103), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1079), .B1(new_n598), .B2(new_n1103), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1048), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n981), .A2(new_n984), .A3(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1043), .A2(G171), .A3(new_n1005), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI211_X1 g690(.A(G1976), .B(G288), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1031), .B1(new_n1116), .B2(new_n1028), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1014), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1042), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n971), .A2(G286), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1043), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1014), .A2(new_n1042), .A3(new_n1122), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(new_n1120), .C1(new_n1013), .C2(new_n1010), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1115), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n947), .B1(new_n1110), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n944), .B(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n931), .A2(G1986), .A3(G290), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT48), .Z(new_n1132));
  NOR2_X1   g707(.A1(new_n698), .A2(new_n938), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n937), .A2(new_n943), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G2067), .B2(new_n761), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1130), .A2(new_n1132), .B1(new_n932), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n942), .B(KEYINPUT46), .Z(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n934), .A2(new_n742), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n932), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT47), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1143), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT47), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n1141), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1136), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1128), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g725(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1152));
  XNOR2_X1  g726(.A(new_n1152), .B(KEYINPUT127), .ZN(new_n1153));
  NOR2_X1   g727(.A1(G229), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n850), .A3(new_n1154), .ZN(G225));
  INV_X1    g729(.A(G225), .ZN(G308));
endmodule


