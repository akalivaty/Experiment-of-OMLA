//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT10), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AND4_X1   g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n193), .C2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G128), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n195), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n202), .A2(new_n203), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n199), .A2(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT79), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n201), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n190), .A3(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n215), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT80), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n189), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n196), .A2(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n201), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n221), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n228), .A3(KEYINPUT10), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n233), .A3(G101), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G128), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n220), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n220), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n201), .A2(new_n242), .A3(KEYINPUT65), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n229), .B1(new_n235), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n255), .A4(new_n252), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n225), .A2(new_n246), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  INV_X1    g073(.A(G227), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G953), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n223), .A2(new_n228), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n216), .B2(new_n224), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(new_n256), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n203), .B1(new_n202), .B2(new_n215), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n222), .A2(KEYINPUT80), .A3(new_n223), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n270), .B1(new_n273), .B2(new_n257), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n272), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n257), .B1(new_n276), .B2(new_n266), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n225), .A2(new_n246), .A3(KEYINPUT83), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT10), .B1(new_n271), .B2(new_n272), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(new_n245), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n285), .A3(new_n268), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n263), .B1(new_n286), .B2(new_n258), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(new_n274), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT81), .B1(new_n277), .B2(KEYINPUT12), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n258), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n262), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n264), .A2(KEYINPUT82), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n258), .A2(new_n294), .A3(new_n263), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n295), .A3(new_n286), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(G469), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(G469), .A2(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  OAI21_X1  g114(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G214), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n193), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT18), .A2(G131), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n306), .B2(new_n308), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT76), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n191), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n204), .ZN(new_n326));
  INV_X1    g140(.A(new_n308), .ZN(new_n327));
  AOI21_X1  g141(.A(G143), .B1(new_n307), .B2(G214), .ZN(new_n328));
  OAI21_X1  g142(.A(G131), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n306), .A2(new_n255), .A3(new_n308), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT17), .B(G131), .C1(new_n327), .C2(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(KEYINPUT16), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT75), .A3(G146), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT16), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G146), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n338), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n324), .B(new_n326), .C1(new_n334), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n342), .B2(new_n341), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n349), .A2(new_n332), .A3(new_n338), .A4(new_n333), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n326), .B1(new_n350), .B2(new_n324), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n188), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G475), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n329), .A2(new_n331), .B1(G146), .B2(new_n337), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n318), .A2(new_n355), .A3(new_n320), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n317), .A2(KEYINPUT19), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n191), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n354), .A2(new_n358), .B1(new_n312), .B2(new_n323), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n347), .B1(new_n326), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n360), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n353), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n193), .A2(G128), .ZN(new_n367));
  INV_X1    g181(.A(G128), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G143), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT90), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT90), .B1(new_n367), .B2(new_n369), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n371), .A2(new_n248), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G134), .B1(new_n376), .B2(new_n370), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT91), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n379), .A2(KEYINPUT87), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(KEYINPUT87), .ZN(new_n381));
  OAI21_X1  g195(.A(G116), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT88), .B1(new_n379), .B2(G116), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  INV_X1    g198(.A(G116), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G122), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT92), .A4(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n383), .A2(new_n386), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n382), .B(new_n388), .C1(new_n389), .C2(new_n387), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT92), .B1(new_n389), .B2(new_n387), .ZN(new_n391));
  OAI21_X1  g205(.A(G107), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n383), .A2(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n382), .A2(new_n207), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n248), .B1(new_n371), .B2(new_n372), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n376), .A2(G134), .A3(new_n370), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n378), .A2(new_n392), .A3(new_n394), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n382), .A2(new_n393), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n394), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n367), .B2(new_n403), .ZN(new_n405));
  AOI211_X1 g219(.A(KEYINPUT89), .B(KEYINPUT13), .C1(new_n193), .C2(G128), .ZN(new_n406));
  OAI221_X1 g220(.A(new_n369), .B1(new_n403), .B2(new_n367), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G134), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n408), .A3(new_n395), .ZN(new_n409));
  INV_X1    g223(.A(G217), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n300), .A2(new_n410), .A3(G953), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n399), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n399), .B2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n188), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G478), .ZN(new_n415));
  NOR2_X1   g229(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n188), .B(new_n421), .C1(new_n412), .C2(new_n413), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n366), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G210), .B1(G237), .B2(G902), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G119), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n426));
  INV_X1    g240(.A(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G116), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n426), .B(G113), .C1(KEYINPUT5), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT2), .A2(G113), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT67), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT2), .A3(G113), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n435));
  INV_X1    g249(.A(G113), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n437), .A3(new_n425), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n223), .A2(new_n429), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n434), .A2(new_n437), .A3(new_n425), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n425), .B1(new_n434), .B2(new_n437), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n439), .B(new_n440), .C1(new_n235), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n228), .A2(new_n315), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n238), .A2(new_n243), .A3(G125), .A4(new_n240), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT85), .B(G224), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(KEYINPUT7), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(KEYINPUT7), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n444), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n440), .B(KEYINPUT8), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n429), .A2(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n215), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n439), .B1(new_n235), .B2(new_n443), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n447), .B(new_n450), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n463), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n444), .A2(KEYINPUT6), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n424), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n424), .A3(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(G234), .A2(G237), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(G952), .A3(new_n304), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(G898), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(G902), .A3(G953), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT94), .Z(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n302), .A2(new_n423), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n410), .B1(G234), .B2(new_n188), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n368), .A2(G119), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n368), .A2(KEYINPUT73), .A3(G119), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n368), .A3(G119), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT74), .B1(new_n427), .B2(G128), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n489), .B(new_n490), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT23), .B1(new_n368), .B2(G119), .ZN(new_n496));
  AND2_X1   g310(.A1(KEYINPUT23), .A2(G119), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n496), .A2(new_n487), .B1(new_n368), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G110), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n494), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n321), .A2(new_n341), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n494), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n346), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n304), .A2(G221), .A3(G234), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT77), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT22), .B(G137), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n507), .B(new_n508), .Z(new_n511));
  AOI21_X1  g325(.A(new_n503), .B1(new_n349), .B2(new_n338), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n500), .A2(new_n501), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n514), .A3(new_n188), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n486), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n510), .ZN(new_n520));
  INV_X1    g334(.A(new_n514), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n485), .A2(G902), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n519), .A2(KEYINPUT78), .A3(new_n524), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n248), .A2(G137), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n250), .A2(G134), .ZN(new_n532));
  OAI21_X1  g346(.A(G131), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n196), .A2(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n256), .B(new_n533), .C1(new_n195), .C2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n443), .B(new_n535), .C1(new_n257), .C2(new_n244), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n535), .B1(new_n257), .B2(new_n244), .ZN(new_n540));
  INV_X1    g354(.A(new_n443), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n536), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n543), .B2(KEYINPUT28), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT69), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n307), .A2(G210), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n546), .A2(new_n547), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n256), .A2(new_n533), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n256), .A2(new_n533), .A3(KEYINPUT66), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n228), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n268), .A2(new_n238), .A3(new_n240), .A4(new_n243), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n443), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n536), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT28), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n557), .B1(new_n566), .B2(new_n538), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n558), .A2(new_n559), .B1(new_n227), .B2(new_n221), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n561), .A2(new_n568), .B1(new_n569), .B2(new_n268), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n536), .B1(new_n570), .B2(new_n443), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT70), .B1(new_n571), .B2(KEYINPUT28), .ZN(new_n572));
  INV_X1    g386(.A(new_n555), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(KEYINPUT30), .A3(new_n535), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n541), .B(new_n575), .C1(new_n570), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n536), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n573), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n188), .B(new_n556), .C1(new_n574), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n566), .A2(new_n557), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n539), .B1(new_n571), .B2(KEYINPUT28), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n557), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n578), .A2(new_n555), .A3(new_n536), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT31), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n578), .A2(new_n555), .A3(KEYINPUT31), .A4(new_n536), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n588), .A2(new_n573), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n585), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n591), .A2(new_n592), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n573), .B1(new_n567), .B2(new_n572), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT72), .A3(new_n597), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n584), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT71), .B1(new_n593), .B2(new_n595), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n602), .A2(new_n606), .A3(new_n594), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n596), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n530), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n484), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n209), .ZN(G3));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n607), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n614));
  INV_X1    g428(.A(G472), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(KEYINPUT95), .B(G472), .C1(new_n593), .C2(G902), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n299), .A2(new_n301), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(KEYINPUT96), .A3(new_n619), .A4(new_n529), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n606), .B1(new_n602), .B2(new_n594), .ZN(new_n623));
  AOI211_X1 g437(.A(KEYINPUT71), .B(new_n595), .C1(new_n600), .C2(new_n601), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n529), .A2(new_n299), .A3(new_n301), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n475), .B1(new_n473), .B2(KEYINPUT97), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n462), .A2(new_n424), .A3(new_n470), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n471), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n632), .B2(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n482), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n415), .A2(new_n188), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n399), .A2(new_n409), .ZN(new_n636));
  INV_X1    g450(.A(new_n411), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n399), .A2(new_n409), .A3(new_n411), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n635), .B1(new_n640), .B2(new_n415), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT33), .B1(new_n412), .B2(new_n413), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n638), .A2(new_n643), .A3(new_n639), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n644), .A3(G478), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n365), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n634), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n629), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT98), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI211_X1 g466(.A(KEYINPUT99), .B(new_n361), .C1(new_n360), .C2(new_n362), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n363), .A2(new_n364), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(KEYINPUT99), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n420), .A2(new_n422), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n353), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n634), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n629), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT100), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n502), .A2(new_n505), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n523), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n519), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n622), .A2(new_n625), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n484), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT37), .B(G110), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  AND3_X1   g487(.A1(new_n299), .A2(new_n301), .A3(new_n633), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT72), .B1(new_n602), .B2(new_n597), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n585), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n608), .A3(new_n584), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n480), .A2(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n477), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n657), .A2(new_n668), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n674), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NAND2_X1  g498(.A1(new_n573), .A2(new_n543), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n589), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n677), .A2(new_n608), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n669), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n680), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n619), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n619), .A2(new_n694), .A3(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n632), .B(KEYINPUT38), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n656), .A2(new_n365), .ZN(new_n697));
  INV_X1    g511(.A(new_n475), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n690), .A2(new_n693), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  NAND4_X1  g515(.A1(new_n641), .A2(new_n365), .A3(new_n645), .A4(new_n680), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n668), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n674), .A2(new_n678), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  OAI21_X1  g519(.A(new_n188), .B1(new_n281), .B2(new_n287), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n301), .A3(new_n288), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(KEYINPUT101), .A3(new_n301), .A4(new_n288), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n609), .A2(new_n648), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT102), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n712), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n609), .A2(new_n658), .A3(new_n710), .A4(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  INV_X1    g531(.A(KEYINPUT97), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n698), .B1(new_n631), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n474), .B2(new_n718), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n482), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n423), .A2(new_n722), .A3(new_n668), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n678), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NOR2_X1   g539(.A1(new_n634), .A2(new_n697), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n593), .B2(G902), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n600), .B1(new_n555), .B2(new_n544), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n594), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n544), .A2(new_n555), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n591), .B2(new_n592), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n732), .B2(new_n595), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n525), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n726), .A2(new_n736), .A3(new_n710), .A4(new_n711), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  INV_X1    g552(.A(new_n702), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n669), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n721), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n633), .A2(new_n707), .A3(new_n301), .A4(new_n288), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n703), .A2(new_n727), .A3(new_n729), .A4(new_n733), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT104), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND2_X1  g562(.A1(new_n602), .A2(new_n597), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n596), .B1(new_n593), .B2(new_n595), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n584), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n525), .B(new_n739), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n631), .A2(new_n471), .A3(new_n698), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n299), .A2(new_n301), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT42), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n702), .A2(KEYINPUT42), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n609), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n255), .ZN(G33));
  NOR2_X1   g576(.A1(new_n657), .A2(new_n681), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n756), .A2(new_n678), .A3(new_n529), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n646), .A2(new_n366), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n646), .A2(new_n768), .A3(new_n366), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n669), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n618), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n292), .A2(new_n296), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n292), .A2(KEYINPUT45), .A3(new_n296), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n298), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  INV_X1    g593(.A(new_n301), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n288), .A2(new_n298), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n780), .B1(new_n782), .B2(new_n777), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n691), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(KEYINPUT106), .A3(new_n755), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT106), .B1(new_n786), .B2(new_n755), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT107), .B(G137), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G39));
  NAND2_X1  g605(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n779), .A2(new_n783), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n678), .A2(new_n529), .A3(new_n702), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n708), .A2(new_n477), .A3(new_n796), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n689), .A2(new_n529), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n646), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n366), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n770), .A2(new_n734), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n801), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n767), .A2(new_n769), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n477), .ZN(new_n809));
  INV_X1    g623(.A(new_n708), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n696), .A2(new_n698), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n736), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n812), .B2(KEYINPUT114), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n807), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n809), .A2(new_n736), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n707), .A2(new_n288), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT109), .Z(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n301), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n755), .B(new_n821), .C1(new_n795), .C2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n818), .B2(new_n819), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n800), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n633), .A3(new_n810), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT117), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n751), .A2(new_n753), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n735), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n810), .A3(new_n755), .A4(new_n809), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT48), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n304), .A2(G952), .ZN(new_n834));
  INV_X1    g648(.A(new_n647), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n802), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n807), .A2(new_n813), .A3(new_n814), .A4(new_n800), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n825), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n827), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n674), .B(new_n678), .C1(new_n682), .C2(new_n703), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n720), .A2(new_n681), .A3(new_n697), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n688), .A2(new_n619), .A3(new_n842), .A4(new_n668), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n742), .B1(new_n721), .B2(new_n741), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT104), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n841), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n712), .A2(new_n716), .A3(new_n724), .A4(new_n737), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n423), .B1(new_n646), .B2(new_n366), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n483), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n620), .A2(new_n628), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n484), .B1(new_n609), .B2(new_n670), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n681), .B1(new_n352), .B2(G475), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n420), .A2(new_n422), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n655), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT110), .B1(new_n863), .B2(new_n796), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n755), .A2(new_n865), .A3(new_n655), .A4(new_n862), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n668), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n678), .A3(new_n619), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n756), .A2(new_n741), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n764), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT111), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n764), .A2(new_n868), .A3(new_n872), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n761), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n852), .A2(new_n853), .A3(new_n860), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n846), .A2(new_n850), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n747), .A2(KEYINPUT52), .A3(new_n841), .A4(new_n843), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(new_n878), .A3(new_n860), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT53), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n880), .A3(KEYINPUT54), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n854), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n737), .A2(new_n724), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT113), .A3(new_n712), .A4(new_n716), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n859), .A2(new_n853), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n852), .A2(new_n874), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n879), .A2(new_n853), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n881), .B1(new_n890), .B2(KEYINPUT54), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n840), .A2(new_n891), .B1(G952), .B2(G953), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n894));
  INV_X1    g708(.A(new_n766), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n735), .A2(new_n780), .A3(new_n698), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n689), .A2(new_n696), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n188), .B1(new_n888), .B2(new_n889), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n467), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n304), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n901), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n906), .A2(new_n911), .ZN(G51));
  XOR2_X1   g726(.A(new_n298), .B(KEYINPUT57), .Z(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n888), .A2(new_n889), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n888), .B2(new_n889), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT119), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n281), .A2(new_n287), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n913), .C1(new_n915), .C2(new_n916), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n900), .A2(G469), .A3(new_n776), .A4(new_n775), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n907), .B1(new_n922), .B2(new_n923), .ZN(G54));
  AND2_X1   g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n900), .A2(new_n360), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n360), .B1(new_n900), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n907), .ZN(G60));
  NAND2_X1  g742(.A1(new_n642), .A2(new_n644), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n635), .B(KEYINPUT59), .Z(new_n930));
  OAI211_X1 g744(.A(new_n929), .B(new_n930), .C1(new_n915), .C2(new_n916), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n908), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n891), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G63));
  XNOR2_X1  g748(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n888), .B2(new_n889), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n520), .A2(new_n521), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n908), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n937), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n890), .A2(new_n665), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT120), .B(new_n935), .C1(new_n940), .C2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n942), .B(new_n908), .C1(new_n939), .C2(new_n938), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n935), .B1(new_n946), .B2(KEYINPUT120), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n448), .B2(new_n478), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n860), .B2(G953), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n903), .B1(G898), .B2(new_n304), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(G900), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n260), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT123), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n758), .A2(new_n760), .A3(new_n764), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n633), .A2(new_n365), .A3(new_n656), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n784), .A2(new_n735), .A3(new_n830), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n747), .A2(new_n841), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n798), .A2(new_n789), .A3(new_n960), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n959), .B1(new_n965), .B2(new_n304), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT124), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT124), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n575), .B1(new_n570), .B2(new_n577), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n356), .A2(new_n357), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n700), .A2(new_n747), .A3(new_n841), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n700), .A2(new_n976), .A3(new_n747), .A4(new_n841), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n798), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n855), .A2(new_n796), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n609), .A2(new_n619), .A3(new_n691), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n789), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n971), .A2(G953), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n973), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n956), .B1(new_n972), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n968), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n971), .B1(new_n966), .B2(KEYINPUT124), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n956), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n985), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n860), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n965), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n579), .B(KEYINPUT126), .Z(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n573), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n907), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n573), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n978), .A2(new_n981), .A3(new_n993), .ZN(new_n999));
  INV_X1    g813(.A(new_n992), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n580), .B2(new_n589), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n875), .A2(new_n880), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT127), .Z(G57));
endmodule


