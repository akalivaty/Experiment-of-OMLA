//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113;
  OR2_X1    g000(.A1(KEYINPUT74), .A2(G125), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT74), .A2(G125), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n192), .B2(G143), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .A4(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n191), .B1(new_n195), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n194), .B2(G143), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n194), .B2(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n205), .B2(new_n190), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n189), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(new_n199), .A3(G143), .ZN(new_n209));
  INV_X1    g023(.A(new_n193), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n197), .A2(new_n199), .A3(new_n196), .A4(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT0), .B(G128), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n198), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n218), .B2(new_n202), .ZN(new_n219));
  INV_X1    g033(.A(new_n189), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n213), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G224), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G953), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n222), .A2(new_n224), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G119), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT70), .A3(G116), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n232), .B2(G116), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(KEYINPUT71), .A3(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT86), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(new_n236), .A3(new_n237), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G113), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n230), .A2(G119), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n239), .A2(new_n241), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g068(.A(G107), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G104), .ZN(new_n256));
  INV_X1    g070(.A(G104), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G107), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT3), .B1(new_n257), .B2(G107), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n257), .C2(G107), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G101), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  XNOR2_X1  g080(.A(G104), .B(G107), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n265), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(G104), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n258), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT83), .A3(G101), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n264), .A2(new_n265), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT4), .B1(new_n264), .B2(new_n265), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n257), .A2(KEYINPUT3), .A3(G107), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n255), .A2(G104), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT82), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g092(.A(new_n263), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n265), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n240), .B1(new_n234), .B2(new_n238), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n241), .A2(new_n242), .A3(new_n236), .A4(new_n237), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G101), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n273), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G122), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n262), .A2(new_n263), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n265), .B1(new_n297), .B2(new_n277), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n298), .A2(new_n287), .B1(new_n283), .B2(new_n284), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n286), .A2(G101), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT4), .A3(new_n280), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n299), .A2(new_n301), .B1(new_n253), .B2(new_n272), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n296), .B1(new_n302), .B2(new_n291), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n295), .B1(new_n303), .B2(KEYINPUT87), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n302), .A2(new_n291), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n228), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT7), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT90), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n224), .B1(new_n222), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n291), .B(KEYINPUT8), .Z(new_n312));
  NAND2_X1  g126(.A1(new_n268), .A2(new_n271), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n280), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n253), .B2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n236), .A4(new_n237), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n239), .A2(new_n241), .B1(new_n316), .B2(new_n252), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT89), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n272), .B1(new_n317), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n322));
  OAI221_X1 g136(.A(new_n322), .B1(new_n223), .B2(G953), .C1(new_n207), .C2(new_n221), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n311), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n273), .B(new_n291), .C1(new_n282), .C2(new_n289), .ZN(new_n325));
  INV_X1    g139(.A(new_n222), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(KEYINPUT7), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(G902), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G210), .B1(G237), .B2(G902), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n308), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n302), .A2(new_n291), .A3(new_n293), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n325), .A2(new_n306), .A3(KEYINPUT6), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n290), .A2(new_n292), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n227), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G902), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n311), .A2(new_n321), .A3(new_n323), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n327), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n332), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n343), .A3(KEYINPUT91), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n339), .A2(new_n342), .A3(new_n332), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT91), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(G214), .B1(G237), .B2(G902), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(G952), .ZN(new_n353));
  INV_X1    g167(.A(G234), .ZN(new_n354));
  INV_X1    g168(.A(G237), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT73), .B(G902), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n352), .B(new_n358), .C1(G234), .C2(G237), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT21), .B(G898), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n361), .B(KEYINPUT103), .Z(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n352), .A3(G214), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(G143), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT17), .A3(G131), .ZN(new_n368));
  INV_X1    g182(.A(G131), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n366), .B(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n370), .B2(KEYINPUT17), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT16), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT74), .A2(G125), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT74), .A2(G125), .ZN(new_n374));
  OAI21_X1  g188(.A(G140), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(G125), .A2(G140), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n187), .B2(new_n188), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT76), .B(new_n192), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(new_n376), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n384), .B2(G146), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT75), .B1(new_n384), .B2(G146), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n387));
  NOR4_X1   g201(.A1(new_n377), .A2(new_n387), .A3(new_n192), .A4(new_n380), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n381), .B(new_n385), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT95), .ZN(new_n390));
  INV_X1    g204(.A(new_n380), .ZN(new_n391));
  NOR2_X1   g205(.A1(G125), .A2(G140), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n189), .B2(G140), .ZN(new_n393));
  OAI211_X1 g207(.A(G146), .B(new_n391), .C1(new_n393), .C2(new_n372), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n384), .A2(KEYINPUT75), .A3(G146), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n381), .A4(new_n385), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n371), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(G125), .A2(G140), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n376), .A2(KEYINPUT77), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n403));
  AND2_X1   g217(.A1(G125), .A2(G140), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n392), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n194), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(KEYINPUT78), .A3(new_n194), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n409), .A2(new_n410), .B1(G146), .B2(new_n393), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT18), .A2(G131), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n366), .B(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n257), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n416), .B(KEYINPUT94), .Z(new_n417));
  NOR3_X1   g231(.A1(new_n400), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT19), .B1(new_n402), .B2(new_n405), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(KEYINPUT19), .B2(new_n393), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n194), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT93), .B1(new_n420), .B2(new_n194), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n394), .B(new_n370), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n414), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n416), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n363), .B(new_n364), .C1(new_n418), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n364), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n390), .A2(new_n399), .ZN(new_n430));
  INV_X1    g244(.A(new_n371), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n417), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n427), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n437));
  OAI21_X1  g251(.A(new_n428), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n416), .B1(new_n432), .B2(new_n426), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n340), .B1(new_n439), .B2(new_n418), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G475), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n442));
  INV_X1    g256(.A(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G116), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n230), .A2(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(G107), .B(new_n442), .C1(new_n446), .C2(KEYINPUT14), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT100), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n190), .B2(G143), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n215), .A2(KEYINPUT97), .A3(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n190), .A2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G134), .ZN(new_n456));
  INV_X1    g270(.A(G134), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G116), .B(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT96), .ZN(new_n463));
  AOI21_X1  g277(.A(G107), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n447), .A2(new_n448), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n449), .A2(new_n459), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n458), .A2(KEYINPUT99), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT99), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n453), .A2(new_n469), .A3(new_n457), .A4(new_n454), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n461), .A2(new_n463), .A3(G107), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n468), .B(new_n470), .C1(new_n471), .C2(new_n464), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT98), .A4(KEYINPUT13), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(new_n454), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n453), .B2(new_n473), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n457), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n467), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT9), .B(G234), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n481), .A2(new_n482), .A3(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT101), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n467), .B(new_n486), .C1(new_n472), .C2(new_n479), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(KEYINPUT102), .A3(new_n487), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n480), .A2(KEYINPUT102), .A3(new_n484), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n358), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n490), .B(new_n493), .ZN(new_n494));
  AND4_X1   g308(.A1(new_n362), .A2(new_n438), .A3(new_n441), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n481), .B2(G902), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT81), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(new_n340), .ZN(new_n499));
  INV_X1    g313(.A(new_n358), .ZN(new_n500));
  XNOR2_X1  g314(.A(G110), .B(G140), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n352), .A2(G227), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT11), .B1(new_n457), .B2(G137), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT11), .ZN(new_n505));
  INV_X1    g319(.A(G137), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(G134), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n504), .A2(new_n507), .B1(new_n457), .B2(G137), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n211), .A2(new_n212), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n201), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n272), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT10), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT84), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n208), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n195), .B2(new_n200), .ZN(new_n522));
  INV_X1    g336(.A(new_n214), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n203), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n288), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n515), .B1(new_n201), .B2(new_n206), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n525), .A2(new_n301), .B1(new_n272), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n509), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n518), .B1(new_n514), .B2(new_n515), .ZN(new_n529));
  AOI211_X1 g343(.A(KEYINPUT84), .B(KEYINPUT10), .C1(new_n513), .C2(new_n272), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n527), .B(new_n509), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n503), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n314), .A2(new_n201), .A3(new_n206), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n514), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n504), .A2(new_n507), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n457), .A2(G137), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G131), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n508), .A2(new_n369), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n509), .B1(new_n514), .B2(new_n534), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT12), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n503), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n531), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n500), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n499), .B1(new_n550), .B2(new_n498), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n531), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT85), .B1(new_n547), .B2(new_n531), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n503), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n531), .A2(new_n548), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n528), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(G469), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n497), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n351), .A2(new_n495), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n522), .A2(new_n524), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT67), .B1(new_n561), .B2(new_n509), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n213), .A2(new_n219), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT67), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n541), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n201), .A2(new_n206), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT69), .B1(new_n506), .B2(G134), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n457), .B2(G137), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n457), .A3(G137), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n506), .A2(KEYINPUT68), .A3(G134), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n567), .A2(new_n569), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G131), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n540), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n562), .A2(new_n565), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n581), .A2(G128), .B1(new_n218), .B2(new_n202), .ZN(new_n582));
  INV_X1    g396(.A(new_n191), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n211), .B2(new_n212), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n540), .A2(new_n574), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n541), .A2(new_n522), .A3(new_n524), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n566), .A2(KEYINPUT72), .A3(new_n575), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n587), .A2(KEYINPUT30), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n285), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n285), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(new_n592), .A3(new_n588), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n355), .A2(new_n352), .A3(G210), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT27), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT26), .B(G101), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n593), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n588), .A2(KEYINPUT67), .B1(new_n566), .B2(new_n575), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n592), .B1(new_n602), .B2(new_n565), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT28), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n576), .A2(new_n592), .A3(new_n588), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT28), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n607), .A3(new_n598), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT29), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n607), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n285), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n593), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(KEYINPUT28), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n599), .A2(new_n609), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n500), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n577), .A2(new_n285), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n606), .B1(new_n620), .B2(new_n593), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n599), .B1(new_n621), .B2(new_n611), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n593), .A2(new_n598), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n591), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT31), .B1(new_n591), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n627));
  NOR2_X1   g441(.A1(G472), .A2(G902), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n619), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT22), .B(G137), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT23), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n232), .B2(G128), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n636), .B(new_n637), .C1(G119), .C2(new_n190), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G110), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT24), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(G119), .B(G128), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n391), .B1(new_n393), .B2(new_n372), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT76), .B1(new_n644), .B2(new_n192), .ZN(new_n645));
  INV_X1    g459(.A(new_n381), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n647), .B2(new_n397), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT79), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n406), .A2(KEYINPUT78), .A3(new_n194), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT78), .B1(new_n406), .B2(new_n194), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI22_X1  g466(.A1(new_n638), .A2(G110), .B1(new_n641), .B2(new_n640), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n394), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n409), .A2(new_n410), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n656), .A2(KEYINPUT79), .A3(new_n394), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n634), .B1(new_n648), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n643), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n389), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n634), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(new_n655), .A3(new_n657), .A4(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n358), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT25), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n659), .A2(new_n663), .A3(KEYINPUT25), .A4(new_n358), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n482), .B1(new_n358), .B2(G234), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(G902), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT80), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n659), .A2(new_n672), .A3(new_n663), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n672), .B1(new_n659), .B2(new_n663), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n631), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n265), .ZN(G3));
  NAND2_X1  g494(.A1(new_n591), .A2(new_n623), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n591), .A2(new_n623), .A3(KEYINPUT31), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n604), .A2(new_n607), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n683), .A2(new_n684), .B1(new_n685), .B2(new_n599), .ZN(new_n686));
  INV_X1    g500(.A(new_n628), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n626), .B2(new_n358), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n559), .A2(new_n677), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n330), .B1(new_n308), .B2(new_n329), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n349), .B1(new_n694), .B2(new_n345), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n331), .A2(new_n343), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n349), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n362), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT33), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n488), .A2(new_n489), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n485), .A2(KEYINPUT33), .A3(new_n487), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n500), .A2(new_n491), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n490), .A2(new_n491), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n438), .B2(new_n441), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n693), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT34), .B(G104), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G6));
  INV_X1    g528(.A(new_n437), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n414), .B1(new_n430), .B2(new_n431), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n427), .B1(new_n716), .B2(new_n433), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n717), .B2(new_n429), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n364), .B(new_n437), .C1(new_n418), .C2(new_n427), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n494), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n441), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n362), .A3(new_n699), .A4(new_n696), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n692), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT35), .B(G107), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G9));
  INV_X1    g540(.A(new_n669), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n666), .B2(new_n667), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n648), .A2(new_n658), .B1(KEYINPUT36), .B2(new_n634), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n634), .A2(KEYINPUT36), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n661), .A2(new_n655), .A3(new_n657), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n671), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT105), .A4(new_n671), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n688), .A2(new_n690), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n351), .A3(new_n495), .A4(new_n559), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT37), .B(G110), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G12));
  OAI21_X1  g555(.A(KEYINPUT32), .B1(new_n686), .B2(new_n687), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n737), .B1(new_n744), .B2(new_n619), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n350), .B1(new_n331), .B2(new_n343), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT104), .ZN(new_n747));
  INV_X1    g561(.A(G900), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n357), .B1(new_n359), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n720), .A2(new_n441), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n494), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n745), .A2(new_n559), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G128), .ZN(G30));
  XOR2_X1   g568(.A(new_n749), .B(KEYINPUT39), .Z(new_n755));
  NAND2_X1  g569(.A1(new_n559), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT40), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n348), .B(KEYINPUT38), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n340), .B1(new_n614), .B2(new_n598), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n599), .B1(new_n591), .B2(new_n593), .ZN(new_n760));
  OAI21_X1  g574(.A(G472), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n494), .B1(new_n438), .B2(new_n441), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n349), .A3(new_n737), .A4(new_n763), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n757), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G143), .ZN(G45));
  AOI211_X1 g580(.A(new_n749), .B(new_n708), .C1(new_n438), .C2(new_n441), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n745), .A2(new_n559), .A3(new_n747), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G146), .ZN(G48));
  NAND3_X1  g583(.A1(new_n747), .A2(new_n362), .A3(new_n709), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n527), .B1(new_n530), .B2(new_n529), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n541), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n531), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n272), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n288), .A2(new_n522), .A3(new_n524), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n282), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n517), .B2(new_n519), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n503), .B1(new_n777), .B2(new_n509), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n773), .A2(new_n503), .B1(new_n778), .B2(new_n547), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n779), .B2(new_n500), .ZN(new_n780));
  INV_X1    g594(.A(new_n549), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n548), .B1(new_n772), .B2(new_n531), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n498), .B(new_n358), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(KEYINPUT106), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n785), .B(G469), .C1(new_n779), .C2(new_n500), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n631), .A3(new_n677), .A4(new_n496), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n770), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT41), .B(G113), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G15));
  NAND3_X1  g605(.A1(new_n720), .A2(new_n721), .A3(new_n441), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n700), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n676), .B1(new_n744), .B2(new_n619), .ZN(new_n795));
  INV_X1    g609(.A(new_n496), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n784), .B2(new_n786), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT107), .B1(new_n788), .B2(new_n723), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G116), .ZN(G18));
  NAND2_X1  g615(.A1(new_n747), .A2(new_n797), .ZN(new_n802));
  INV_X1    g616(.A(new_n736), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n670), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n631), .A2(new_n495), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n232), .ZN(G21));
  NAND2_X1  g621(.A1(new_n683), .A2(new_n684), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n606), .B1(new_n613), .B2(new_n593), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n599), .B1(new_n809), .B2(new_n611), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n687), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n676), .A2(new_n690), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n797), .A2(new_n362), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n747), .A2(new_n763), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n443), .ZN(G24));
  NOR3_X1   g630(.A1(new_n690), .A2(new_n737), .A3(new_n811), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n747), .A2(new_n797), .A3(new_n767), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G125), .ZN(G27));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT42), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(KEYINPUT108), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n796), .B1(new_n551), .B2(new_n558), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n350), .B1(new_n344), .B2(new_n347), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n631), .A2(new_n823), .A3(new_n677), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n438), .A2(new_n441), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n707), .A3(new_n750), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n822), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n499), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n558), .A2(new_n829), .A3(new_n783), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n824), .A2(new_n830), .A3(new_n496), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n822), .B1(new_n820), .B2(new_n821), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n795), .A3(new_n767), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n369), .ZN(G33));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n795), .A3(new_n752), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G134), .ZN(G36));
  NOR2_X1   g651(.A1(new_n691), .A2(new_n737), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n438), .A2(new_n441), .A3(new_n707), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT43), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT43), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT44), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n824), .B(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n842), .A2(new_n847), .A3(new_n843), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n842), .B2(new_n843), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT45), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT85), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n545), .B(new_n543), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n532), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n531), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n548), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n851), .B1(new_n856), .B2(new_n556), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n554), .A2(KEYINPUT45), .A3(new_n557), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(G469), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT46), .B1(new_n859), .B2(new_n829), .ZN(new_n860));
  INV_X1    g674(.A(new_n783), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(KEYINPUT46), .A3(new_n829), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n796), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n755), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n864), .B2(new_n755), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n850), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(G137), .ZN(G39));
  OR2_X1    g683(.A1(new_n864), .A2(KEYINPUT47), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(KEYINPUT47), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n348), .A2(new_n349), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n631), .A2(new_n827), .A3(new_n873), .A4(new_n677), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(G140), .ZN(G42));
  XNOR2_X1  g690(.A(new_n787), .B(KEYINPUT49), .ZN(new_n877));
  INV_X1    g691(.A(new_n497), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n677), .A2(new_n349), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n762), .A2(new_n879), .A3(new_n839), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n880), .A3(new_n758), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n787), .A2(new_n497), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n870), .A2(new_n871), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n840), .A2(new_n357), .A3(new_n812), .A4(new_n841), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n845), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n758), .A2(new_n350), .A3(new_n797), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n889), .A2(new_n890), .A3(new_n884), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n889), .B2(new_n884), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n357), .A3(new_n841), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n797), .A2(new_n824), .ZN(new_n895));
  OAI21_X1  g709(.A(G472), .B1(new_n686), .B2(new_n500), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n808), .A2(new_n810), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n628), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n804), .A3(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n677), .A2(new_n357), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n895), .A2(new_n762), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n826), .A2(new_n707), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n888), .A2(new_n893), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n888), .A2(KEYINPUT51), .A3(new_n893), .A4(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n709), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n909), .B(new_n353), .C1(new_n802), .C2(new_n884), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n894), .A2(new_n895), .A3(new_n678), .ZN(new_n911));
  XOR2_X1   g725(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n907), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT119), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n907), .A2(new_n908), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n783), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n533), .A2(new_n549), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n498), .B1(new_n923), .B2(new_n358), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n786), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n496), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n678), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n696), .A2(new_n699), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n631), .A2(new_n495), .A3(new_n804), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n711), .A2(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n739), .B1(new_n560), .B2(new_n678), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n362), .B(new_n496), .C1(new_n925), .C2(new_n926), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n690), .A2(new_n811), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n677), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n696), .A2(new_n763), .A3(new_n699), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n438), .A2(new_n441), .A3(new_n494), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n344), .A2(new_n347), .A3(new_n349), .A4(new_n362), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n707), .B1(new_n438), .B2(new_n441), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n938), .A2(new_n939), .B1(new_n693), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n800), .A2(new_n932), .A3(new_n934), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n827), .A2(new_n899), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT113), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n831), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n936), .A2(new_n709), .A3(new_n804), .A4(new_n750), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n824), .A2(new_n830), .A3(new_n496), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT113), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n856), .A2(new_n498), .A3(new_n556), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n783), .A2(new_n829), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n494), .B(new_n878), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n873), .A3(new_n751), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n949), .A2(new_n952), .B1(new_n745), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(new_n828), .A3(new_n833), .A4(new_n836), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n946), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n728), .A2(new_n736), .A3(new_n749), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n496), .C1(new_n953), .C2(new_n954), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n939), .A2(new_n962), .A3(new_n762), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n753), .A2(new_n768), .A3(new_n963), .A4(new_n818), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT115), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT52), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n753), .A2(new_n818), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(KEYINPUT52), .A3(new_n768), .A4(new_n963), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n965), .A2(new_n967), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT53), .B(new_n959), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT116), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n968), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n974), .B(KEYINPUT53), .C1(new_n959), .C2(new_n975), .ZN(new_n976));
  AND4_X1   g790(.A1(new_n800), .A2(new_n932), .A3(new_n934), .A4(new_n945), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n949), .A2(new_n952), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n956), .A2(new_n745), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n828), .A2(new_n833), .A3(new_n836), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n975), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT53), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT116), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n921), .B(new_n973), .C1(new_n976), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n988));
  OAI22_X1  g802(.A1(new_n770), .A2(new_n788), .B1(new_n802), .B2(new_n805), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n826), .A2(new_n708), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n351), .A2(new_n362), .A3(new_n940), .A4(new_n990), .ZN(new_n991));
  OAI22_X1  g805(.A1(new_n813), .A2(new_n814), .B1(new_n991), .B2(new_n692), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n989), .A2(new_n992), .A3(new_n933), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n982), .A2(new_n800), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT114), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n988), .B(new_n996), .C1(new_n971), .C2(new_n972), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n987), .B1(new_n997), .B2(new_n984), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n986), .B1(new_n998), .B2(new_n921), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n920), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(G952), .A2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n881), .B1(new_n1000), .B2(new_n1001), .ZN(G75));
  OAI21_X1  g816(.A(new_n973), .B1(new_n976), .B2(new_n985), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n500), .A3(new_n332), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT56), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n304), .A2(new_n228), .A3(new_n307), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n339), .ZN(new_n1007));
  XNOR2_X1  g821(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1004), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n352), .A2(G952), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(G51));
  XNOR2_X1  g827(.A(new_n499), .B(KEYINPUT57), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n964), .B(KEYINPUT52), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n984), .B1(new_n994), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n974), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n983), .A2(KEYINPUT116), .A3(new_n984), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n921), .B1(new_n1019), .B2(new_n973), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n982), .A2(new_n993), .A3(KEYINPUT53), .A4(new_n800), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n975), .A2(new_n965), .ZN(new_n1022));
  INV_X1    g836(.A(new_n972), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g838(.A(KEYINPUT54), .B(new_n1024), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1014), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n923), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1003), .A2(new_n500), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n1028), .A2(new_n859), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1012), .B1(new_n1027), .B2(new_n1029), .ZN(G54));
  NAND2_X1  g844(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n717), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1012), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1028), .A2(new_n717), .A3(new_n1031), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1034), .A2(new_n1035), .ZN(G60));
  NAND2_X1  g850(.A1(G478), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT59), .Z(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  AOI22_X1  g853(.A1(new_n999), .A2(new_n1039), .B1(new_n702), .B2(new_n703), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n702), .A2(new_n703), .A3(new_n1039), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1003), .A2(KEYINPUT54), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1042), .B2(new_n986), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1040), .A2(new_n1012), .A3(new_n1043), .ZN(G63));
  XNOR2_X1  g858(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G217), .A2(G902), .ZN(new_n1046));
  XNOR2_X1  g860(.A(new_n1046), .B(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1003), .A2(new_n1048), .ZN(new_n1049));
  OR2_X1    g863(.A1(new_n673), .A2(new_n674), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1012), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n729), .A2(new_n731), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1003), .A2(new_n1053), .A3(new_n1048), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1045), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1024), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1051), .B1(new_n1056), .B2(new_n1047), .ZN(new_n1057));
  AND4_X1   g871(.A1(new_n1033), .A2(new_n1057), .A3(new_n1054), .A4(new_n1045), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1055), .A2(new_n1058), .ZN(G66));
  NAND2_X1  g873(.A1(new_n946), .A2(new_n352), .ZN(new_n1060));
  OAI21_X1  g874(.A(G953), .B1(new_n360), .B2(new_n223), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1060), .A2(KEYINPUT122), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n1062), .B1(KEYINPUT122), .B2(new_n1060), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n335), .B(new_n338), .C1(G898), .C2(new_n352), .ZN(new_n1064));
  XOR2_X1   g878(.A(new_n1063), .B(new_n1064), .Z(G69));
  AOI21_X1  g879(.A(new_n352), .B1(G227), .B2(G900), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n579), .A2(new_n590), .ZN(new_n1067));
  XOR2_X1   g881(.A(new_n1067), .B(new_n420), .Z(new_n1068));
  NAND3_X1  g882(.A1(new_n969), .A2(KEYINPUT123), .A3(new_n768), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n753), .A2(new_n768), .A3(new_n818), .ZN(new_n1070));
  INV_X1    g884(.A(KEYINPUT123), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1073), .A2(new_n765), .ZN(new_n1074));
  INV_X1    g888(.A(KEYINPUT62), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n1073), .A2(KEYINPUT62), .A3(new_n765), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n756), .A2(new_n873), .ZN(new_n1079));
  NAND4_X1  g893(.A1(new_n1079), .A2(new_n795), .A3(new_n940), .A4(new_n990), .ZN(new_n1080));
  NAND4_X1  g894(.A1(new_n1078), .A2(new_n868), .A3(new_n875), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g895(.A(new_n1068), .B1(new_n1081), .B2(new_n352), .ZN(new_n1082));
  OAI211_X1 g896(.A(new_n795), .B(new_n939), .C1(new_n866), .C2(new_n867), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n981), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1084));
  NAND4_X1  g898(.A1(new_n875), .A2(new_n1083), .A3(new_n868), .A4(new_n1084), .ZN(new_n1085));
  NOR2_X1   g899(.A1(new_n1085), .A2(G953), .ZN(new_n1086));
  OAI21_X1  g900(.A(new_n1068), .B1(new_n748), .B2(new_n352), .ZN(new_n1087));
  NOR2_X1   g901(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g902(.A(new_n1066), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g903(.A(new_n1066), .B(KEYINPUT125), .ZN(new_n1090));
  OAI221_X1 g904(.A(new_n1090), .B1(new_n1086), .B2(new_n1087), .C1(new_n1082), .C2(KEYINPUT124), .ZN(new_n1091));
  AND2_X1   g905(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1092));
  OAI21_X1  g906(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(G72));
  NOR2_X1   g907(.A1(new_n594), .A2(new_n598), .ZN(new_n1094));
  XNOR2_X1  g908(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1095));
  NOR2_X1   g909(.A1(new_n689), .A2(new_n340), .ZN(new_n1096));
  XOR2_X1   g910(.A(new_n1095), .B(new_n1096), .Z(new_n1097));
  INV_X1    g911(.A(new_n1097), .ZN(new_n1098));
  OR3_X1    g912(.A1(new_n1094), .A2(new_n760), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g913(.A1(new_n998), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g914(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g915(.A(new_n1097), .B1(new_n1081), .B2(new_n946), .ZN(new_n1102));
  NAND2_X1  g916(.A1(new_n1102), .A2(new_n760), .ZN(new_n1103));
  INV_X1    g917(.A(KEYINPUT127), .ZN(new_n1104));
  OAI21_X1  g918(.A(new_n1097), .B1(new_n1085), .B2(new_n946), .ZN(new_n1105));
  AOI21_X1  g919(.A(new_n1012), .B1(new_n1105), .B2(new_n1094), .ZN(new_n1106));
  NAND4_X1  g920(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g921(.A1(new_n875), .A2(new_n868), .A3(new_n1080), .ZN(new_n1108));
  AOI21_X1  g922(.A(new_n1108), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1109));
  AOI21_X1  g923(.A(new_n1098), .B1(new_n1109), .B2(new_n977), .ZN(new_n1110));
  INV_X1    g924(.A(new_n760), .ZN(new_n1111));
  OAI21_X1  g925(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g926(.A(KEYINPUT127), .B1(new_n1112), .B2(new_n1100), .ZN(new_n1113));
  NAND2_X1  g927(.A1(new_n1107), .A2(new_n1113), .ZN(G57));
endmodule


