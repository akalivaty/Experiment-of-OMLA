//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n628, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT68), .B(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT70), .Z(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n468), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n468), .A2(new_n481), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g064(.A1(G124), .A2(new_n487), .B1(new_n489), .B2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n463), .A2(G2104), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n496), .B2(new_n485), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n468), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT4), .A2(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n469), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n497), .B(new_n501), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n513), .B1(new_n510), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n519), .A2(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT73), .Z(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(new_n526), .A3(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n519), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n533), .B(new_n541), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT7), .Z(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n520), .B2(G89), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n542), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n517), .B2(new_n518), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT76), .B(G52), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n522), .A2(G543), .A3(new_n523), .A4(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n522), .A2(G90), .A3(new_n523), .A4(new_n519), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n518), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT5), .A2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n514), .A2(G81), .A3(new_n519), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n514), .A2(G43), .A3(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT78), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(new_n520), .A2(G91), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  OAI21_X1  g152(.A(G65), .B1(new_n558), .B2(new_n559), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(new_n580), .B2(G651), .ZN(new_n581));
  AOI211_X1 g156(.A(KEYINPUT80), .B(new_n512), .C1(new_n578), .C2(new_n579), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G53), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT9), .B1(new_n524), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n514), .A2(new_n587), .A3(G53), .A4(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(KEYINPUT79), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT79), .B1(new_n586), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(G299));
  XNOR2_X1  g167(.A(new_n555), .B(KEYINPUT81), .ZN(G301));
  NAND3_X1  g168(.A1(new_n514), .A2(G87), .A3(new_n519), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n522), .A2(G49), .A3(G543), .A4(new_n523), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n517), .B2(new_n518), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n523), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n522), .A2(G86), .A3(new_n523), .A4(new_n519), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n520), .A2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n525), .A2(G47), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(new_n512), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n560), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n525), .A2(G54), .B1(new_n612), .B2(G651), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n514), .A2(G92), .A3(new_n519), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n618), .B(G301), .S(G868), .Z(G321));
  XNOR2_X1  g194(.A(G321), .B(KEYINPUT83), .ZN(G284));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n586), .A2(new_n588), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n583), .B1(new_n624), .B2(new_n589), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n621), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n621), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(new_n618), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n474), .A2(new_n471), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  OAI221_X1 g213(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n639));
  INV_X1    g214(.A(G123), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n639), .B1(new_n486), .B2(new_n640), .C1(new_n641), .C2(new_n488), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT86), .B1(new_n651), .B2(KEYINPUT14), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n660), .B(new_n649), .C1(new_n652), .C2(new_n655), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n659), .A2(new_n668), .A3(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G14), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n666), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n674), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(KEYINPUT17), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n676), .B1(new_n675), .B2(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT18), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1981), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT89), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n701), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G20), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT23), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n625), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1956), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2090), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT102), .B(KEYINPUT29), .Z(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(G4), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n628), .B2(new_n707), .ZN(new_n721));
  INV_X1    g296(.A(G1348), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n712), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G128), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n489), .A2(G140), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2067), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n707), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n567), .B2(new_n707), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n723), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT96), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n712), .A2(G32), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n489), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n471), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n738), .B1(new_n747), .B2(new_n712), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT27), .B(G1996), .Z(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT100), .Z(new_n751));
  AND2_X1   g326(.A1(new_n712), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G139), .B2(new_n489), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(new_n469), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT99), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n761), .A2(KEYINPUT99), .A3(new_n762), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n751), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n712), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NOR2_X1   g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n712), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT98), .ZN(new_n773));
  INV_X1    g348(.A(G160), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n712), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n769), .B1(new_n712), .B2(new_n642), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(G164), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G27), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n707), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n707), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n761), .A2(new_n762), .B1(G1961), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT101), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n748), .A2(new_n749), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n775), .A2(new_n776), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n788), .B(new_n789), .C1(G1961), .C2(new_n785), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n783), .B(new_n786), .C1(new_n787), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n707), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n707), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G1966), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n790), .A2(new_n787), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(G1966), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n765), .A2(new_n791), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n719), .A2(new_n737), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n800));
  NAND2_X1  g375(.A1(G288), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n595), .A4(new_n596), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G23), .B(new_n803), .S(G16), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n707), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n707), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G6), .B(G305), .S(G16), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n807), .A2(new_n808), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NOR2_X1   g392(.A1(G16), .A2(G24), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT93), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT92), .B(G1986), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n712), .A2(G25), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT90), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n487), .A2(G119), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n469), .A2(G107), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n489), .A2(G131), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n825), .B1(new_n832), .B2(G29), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n823), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n817), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n799), .B1(new_n839), .B2(new_n840), .ZN(G311));
  INV_X1    g416(.A(new_n799), .ZN(new_n842));
  INV_X1    g417(.A(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(G150));
  NAND2_X1  g420(.A1(new_n628), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n514), .A2(G93), .A3(new_n519), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n514), .A2(G55), .A3(G543), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n848), .B(new_n849), .C1(new_n512), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n566), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  OAI221_X1 g435(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  INV_X1    g437(.A(G142), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n861), .B1(new_n486), .B2(new_n862), .C1(new_n863), .C2(new_n488), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT104), .ZN(new_n865));
  INV_X1    g440(.A(new_n636), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(new_n832), .ZN(new_n870));
  INV_X1    g445(.A(new_n832), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n864), .B(KEYINPUT104), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n636), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n873), .B2(new_n867), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT105), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n832), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n871), .A3(new_n867), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n730), .A2(new_n507), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n730), .A2(new_n507), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n747), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n746), .A3(new_n880), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n760), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n760), .A2(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n883), .B(new_n885), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n875), .A2(new_n879), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n890), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n870), .A2(new_n874), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n877), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n774), .B(new_n642), .ZN(new_n898));
  XNOR2_X1  g473(.A(G162), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g480(.A(G290), .B(G303), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n803), .B(G305), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n853), .B(new_n631), .ZN(new_n911));
  NAND2_X1  g486(.A1(G299), .A2(new_n618), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n625), .A2(new_n628), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT41), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n910), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G868), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n851), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n927), .ZN(G331));
  INV_X1    g504(.A(new_n908), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n545), .A2(new_n542), .ZN(new_n931));
  INV_X1    g506(.A(new_n538), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n536), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n541), .B1(new_n933), .B2(new_n533), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n555), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G301), .B2(G286), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n853), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT81), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n555), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n931), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n540), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n852), .A3(new_n935), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n917), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT41), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n941), .A2(new_n852), .A3(new_n935), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n852), .B1(new_n941), .B2(new_n935), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n914), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n930), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n937), .B(new_n942), .C1(new_n916), .C2(new_n917), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(new_n943), .B2(new_n914), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n908), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n901), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n930), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n955), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n961), .A3(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n957), .A2(new_n961), .A3(KEYINPUT111), .A4(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(new_n956), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n959), .A2(KEYINPUT109), .A3(new_n968), .A4(new_n955), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n967), .C2(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n966), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n507), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n482), .A2(new_n484), .A3(new_n505), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n503), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n500), .B1(new_n982), .B2(new_n468), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n983), .B2(new_n497), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n473), .A2(new_n477), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT120), .B(G1996), .Z(new_n988));
  NAND4_X1  g563(.A1(new_n980), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT121), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n979), .B(G1384), .C1(new_n983), .C2(new_n497), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n507), .B2(new_n977), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(KEYINPUT121), .A3(new_n987), .A4(new_n988), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT58), .B(G1341), .Z(new_n996));
  INV_X1    g571(.A(new_n477), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(G40), .A3(new_n472), .A4(new_n470), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(new_n978), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT59), .A3(new_n567), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n984), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n984), .A2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n987), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n978), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n722), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n998), .A2(new_n978), .ZN(new_n1010));
  INV_X1    g585(.A(G2067), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1009), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1001), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT59), .B1(new_n1000), .B2(new_n567), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  INV_X1    g592(.A(G1956), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n987), .B1(new_n984), .B2(new_n1003), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n501), .B1(new_n506), .B2(new_n502), .ZN(new_n1020));
  INV_X1    g595(.A(new_n497), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1003), .B(new_n977), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1018), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT119), .B(new_n1018), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n625), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n584), .A2(new_n1029), .A3(new_n622), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n992), .A2(new_n993), .A3(new_n998), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1028), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1017), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1032), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1028), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT61), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1022), .A2(KEYINPUT113), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n998), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1007), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(new_n722), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT60), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1052), .A3(new_n628), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1016), .A2(new_n1038), .A3(new_n1043), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1048), .A2(new_n618), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1042), .B1(new_n1055), .B2(new_n1037), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT122), .B(G1961), .Z(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1047), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1033), .A2(new_n780), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1064), .A2(new_n1065), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1061), .B(KEYINPUT123), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(G301), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1062), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1062), .B(new_n986), .C1(KEYINPUT125), .C2(G2078), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n997), .B(new_n1070), .C1(KEYINPUT125), .C2(G2078), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n473), .A2(KEYINPUT124), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n994), .B(new_n1073), .C1(KEYINPUT124), .C2(new_n473), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1061), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n939), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1058), .B1(new_n1068), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n987), .B2(new_n984), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n801), .A2(G1976), .A3(new_n802), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1080), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G305), .A2(G1981), .ZN(new_n1086));
  INV_X1    g661(.A(G1981), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(KEYINPUT49), .A3(new_n1088), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n1080), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT115), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n1092), .A4(new_n1080), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1082), .B(new_n1085), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1971), .B1(new_n994), .B2(new_n987), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1019), .A2(new_n1023), .A3(G2090), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G303), .A2(G8), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT55), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1105));
  INV_X1    g680(.A(G2090), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n987), .A4(new_n1007), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n980), .A2(new_n985), .A3(new_n987), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n811), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1101), .B(KEYINPUT55), .Z(new_n1111));
  AND4_X1   g686(.A1(new_n1104), .A2(new_n1110), .A3(new_n1111), .A4(G8), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1079), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1104), .B1(new_n1113), .B2(new_n1111), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1097), .B(new_n1103), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT116), .B1(new_n1033), .B2(G1966), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  INV_X1    g692(.A(G1966), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1108), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1105), .A2(new_n776), .A3(new_n987), .A4(new_n1007), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1116), .A2(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1046), .A2(KEYINPUT117), .A3(new_n776), .A4(new_n1007), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(G168), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G8), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT51), .ZN(new_n1126));
  AOI21_X1  g701(.A(G168), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n1128));
  OAI211_X1 g703(.A(G8), .B(new_n1124), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1115), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1063), .A2(new_n1062), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1059), .B1(new_n1046), .B2(new_n1007), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1065), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1067), .A2(new_n1134), .A3(new_n1069), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1135), .B2(new_n939), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1066), .A2(KEYINPUT126), .A3(G301), .A4(new_n1067), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1058), .B1(new_n1075), .B2(G171), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1057), .A2(new_n1077), .A3(new_n1130), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n1123), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G286), .A2(new_n1079), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1085), .A2(new_n1082), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1146), .B(new_n1147), .C1(new_n1113), .C2(new_n1111), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT63), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1080), .ZN(new_n1150));
  INV_X1    g725(.A(G288), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1083), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1152), .B2(new_n1088), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1097), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1110), .A2(new_n1111), .A3(G8), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT114), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1113), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1156), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT118), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1161), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1097), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1110), .A2(G8), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1102), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1169), .A2(new_n1097), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1153), .B1(new_n1170), .B2(KEYINPUT63), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1167), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1164), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1128), .B1(new_n1143), .B2(G286), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1125), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1128), .B1(new_n1124), .B2(G8), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT62), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1126), .A2(new_n1129), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1135), .A2(new_n939), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1115), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1178), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1140), .A2(new_n1174), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n980), .A2(new_n998), .ZN(new_n1185));
  INV_X1    g760(.A(new_n834), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n832), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n730), .B(new_n1011), .ZN(new_n1188));
  INV_X1    g763(.A(G1996), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n746), .B(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(G1986), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n819), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT112), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1194), .B2(new_n819), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1185), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1184), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1185), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1201), .B1(new_n1188), .B2(new_n747), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1201), .A2(new_n1203), .A3(G1996), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT46), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1205));
  OR3_X1    g780(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT48), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1196), .A2(KEYINPUT48), .A3(new_n1185), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1210), .B(new_n1211), .C1(new_n1201), .C2(new_n1192), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1191), .A2(new_n1186), .A3(new_n832), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n730), .A2(G2067), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1185), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1216));
  AND4_X1   g791(.A1(new_n1208), .A2(new_n1212), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1200), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g793(.A1(G227), .A2(new_n461), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1220), .B1(new_n671), .B2(new_n672), .ZN(new_n1221));
  OR2_X1    g795(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1222));
  AOI21_X1  g796(.A(G229), .B1(new_n1221), .B2(KEYINPUT127), .ZN(new_n1223));
  AND3_X1   g797(.A1(new_n904), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AND2_X1   g798(.A1(new_n1224), .A2(new_n974), .ZN(G308));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n974), .ZN(G225));
endmodule


