//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n595, new_n596, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(new_n464), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XOR2_X1   g049(.A(KEYINPUT3), .B(G2104), .Z(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G2105), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT66), .ZN(G160));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n468), .A2(new_n470), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(G2105), .A3(new_n466), .ZN(new_n487));
  OAI221_X1 g062(.A(new_n483), .B1(new_n471), .B2(new_n484), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR4_X1   g065(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n490), .A4(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n471), .B2(new_n490), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT67), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n486), .A2(G138), .A3(new_n467), .A4(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n486), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT6), .B(G651), .Z(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(G166));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT68), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G51), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n514), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n505), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT7), .Z(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  AOI22_X1  g100(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n508), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n511), .A2(new_n505), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n527), .B1(G90), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G171));
  NAND2_X1  g107(.A1(new_n528), .A2(G81), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n533), .B1(new_n534), .B2(new_n508), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT69), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT70), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT72), .Z(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n505), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n528), .A2(G91), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n517), .A2(G53), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(G299));
  XOR2_X1   g133(.A(new_n531), .B(KEYINPUT73), .Z(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  NAND2_X1  g135(.A1(new_n517), .A2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n528), .A2(G87), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  AOI22_X1  g139(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n508), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n506), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n511), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G305));
  NAND2_X1  g145(.A1(new_n528), .A2(G85), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT74), .B(G47), .Z(new_n573));
  OAI221_X1 g148(.A(new_n571), .B1(new_n572), .B2(new_n508), .C1(new_n535), .C2(new_n573), .ZN(G290));
  NAND2_X1  g149(.A1(new_n528), .A2(G92), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT10), .Z(new_n576));
  AOI22_X1  g151(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n508), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(G54), .B2(new_n517), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(G868), .ZN(new_n581));
  INV_X1    g156(.A(G301), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(G868), .ZN(G284));
  AOI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(G868), .ZN(G321));
  NAND2_X1  g159(.A1(G286), .A2(G868), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT75), .Z(new_n586));
  OR2_X1    g161(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n552), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n586), .B1(new_n589), .B2(G868), .ZN(G297));
  XOR2_X1   g165(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g166(.A(new_n580), .ZN(new_n592));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G860), .ZN(G148));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G868), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G868), .B2(new_n538), .ZN(G323));
  XNOR2_X1  g172(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g173(.A(new_n487), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G123), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT78), .Z(new_n601));
  NAND2_X1  g176(.A1(new_n472), .A2(G135), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n467), .A2(G111), .ZN(new_n603));
  OAI21_X1  g178(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT79), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(G2096), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(G2096), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT13), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(G2100), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n612), .B2(new_n611), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n613), .A2(G2100), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n609), .A3(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  AOI21_X1  g215(.A(KEYINPUT18), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n636), .A2(new_n637), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XOR2_X1   g222(.A(G1971), .B(G1976), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT19), .ZN(new_n649));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  AND2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  OR3_X1    g232(.A1(new_n649), .A2(new_n652), .A3(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT83), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1981), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  NOR2_X1   g242(.A1(G16), .A2(G24), .ZN(new_n668));
  XNOR2_X1  g243(.A(G290), .B(KEYINPUT85), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n669), .B2(G16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1986), .ZN(new_n671));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G23), .ZN(new_n673));
  INV_X1    g248(.A(G288), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT33), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(G22), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G166), .B2(new_n672), .ZN(new_n680));
  INV_X1    g255(.A(G1971), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n672), .A2(G6), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n569), .B2(new_n672), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n678), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n671), .B1(KEYINPUT34), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G25), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n599), .A2(G119), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n472), .A2(G131), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n689), .B(new_n700), .C1(KEYINPUT34), .C2(new_n688), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT36), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n472), .A2(G141), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n599), .A2(G129), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n708), .A2(new_n709), .B1(G105), .B2(new_n478), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT93), .ZN(new_n712));
  MUX2_X1   g287(.A(G32), .B(new_n712), .S(G29), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT95), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n690), .A2(G26), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT28), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n599), .A2(G128), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n472), .A2(G140), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n467), .A2(G116), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n721), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT89), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2067), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n690), .A2(G27), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT97), .Z(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n690), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G2078), .Z(new_n733));
  NAND4_X1  g308(.A1(new_n717), .A2(new_n718), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n607), .A2(new_n690), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n690), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n690), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT29), .B(G2090), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n690), .B1(new_n740), .B2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n740), .B2(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G160), .B2(G29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G2084), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(G2084), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n735), .A2(new_n739), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n672), .A2(G20), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT23), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n589), .B2(new_n672), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n672), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n538), .B2(new_n672), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT88), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n592), .A2(new_n672), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G4), .B2(new_n672), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n672), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n672), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G33), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT90), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n472), .A2(G139), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  INV_X1    g343(.A(G127), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n475), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n766), .B(new_n768), .C1(new_n771), .C2(new_n467), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n690), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n759), .B(new_n763), .C1(KEYINPUT91), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n672), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n672), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT96), .B(G28), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n782), .B2(KEYINPUT30), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n780), .B(new_n785), .C1(new_n774), .C2(new_n773), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n757), .B2(new_n758), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n776), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n746), .A2(new_n751), .A3(new_n755), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n702), .A2(new_n734), .A3(new_n790), .ZN(G311));
  INV_X1    g366(.A(G311), .ZN(G150));
  AOI22_X1  g367(.A1(new_n517), .A2(G55), .B1(G93), .B2(new_n528), .ZN(new_n793));
  NAND2_X1  g368(.A1(G80), .A2(G543), .ZN(new_n794));
  INV_X1    g369(.A(G67), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n505), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n508), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT101), .B(G860), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT102), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT37), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n538), .A2(new_n800), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n807));
  INV_X1    g382(.A(new_n800), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(new_n537), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n592), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT39), .Z(new_n815));
  OAI21_X1  g390(.A(new_n804), .B1(new_n815), .B2(new_n801), .ZN(G145));
  NAND2_X1  g391(.A1(new_n599), .A2(G130), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n472), .A2(G142), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n467), .A2(G118), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT106), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n611), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n696), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n712), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT105), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n501), .A2(KEYINPUT104), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT104), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n498), .A2(new_n828), .A3(new_n500), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n826), .B1(new_n497), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n491), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT4), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n495), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n498), .A2(new_n828), .A3(new_n500), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n828), .B1(new_n498), .B2(new_n500), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(KEYINPUT105), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n772), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n727), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n825), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G160), .B(KEYINPUT103), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n607), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n843), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT107), .B(G37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g425(.A1(new_n589), .A2(new_n580), .ZN(new_n851));
  NAND2_X1  g426(.A1(G299), .A2(new_n592), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(G299), .A2(KEYINPUT108), .A3(new_n592), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n851), .A2(new_n852), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(KEYINPUT41), .B2(new_n856), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n810), .B(new_n595), .ZN(new_n861));
  MUX2_X1   g436(.A(new_n856), .B(new_n860), .S(new_n861), .Z(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G288), .B(G166), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(new_n569), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n865), .B(new_n866), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n864), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(G868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G868), .B2(new_n808), .ZN(G295));
  OAI21_X1  g447(.A(new_n871), .B1(G868), .B2(new_n808), .ZN(G331));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n810), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(G171), .A2(G168), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n582), .B2(G168), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n810), .B(KEYINPUT109), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n856), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT110), .ZN(new_n884));
  INV_X1    g459(.A(new_n856), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n876), .A2(new_n878), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n879), .A2(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n860), .ZN(new_n892));
  INV_X1    g467(.A(new_n867), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n884), .A2(new_n890), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n860), .A2(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n874), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n857), .A2(KEYINPUT41), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT111), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n879), .A2(new_n882), .A3(new_n858), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n885), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n867), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .A3(new_n848), .A4(new_n894), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n896), .B2(new_n898), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n905), .A2(new_n874), .A3(new_n848), .A4(new_n894), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n913), .ZN(G397));
  OR2_X1    g489(.A1(new_n712), .A2(G1996), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n726), .B(G2067), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n712), .A2(G1996), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n697), .A2(new_n699), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n918), .A2(new_n919), .B1(G2067), .B2(new_n727), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n831), .A2(new_n921), .A3(new_n839), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n473), .A2(new_n479), .A3(G40), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n916), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n930), .B2(new_n712), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n927), .A2(new_n932), .A3(G1996), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n927), .B2(G1996), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT47), .Z(new_n936));
  OR3_X1    g511(.A1(new_n927), .A2(G1986), .A3(G290), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  INV_X1    g515(.A(new_n918), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n697), .A2(new_n699), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n919), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n943), .B2(new_n928), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n929), .B(new_n936), .C1(new_n939), .C2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G290), .B(G1986), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n928), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n950));
  OAI22_X1  g525(.A1(G166), .A2(new_n949), .B1(KEYINPUT113), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(KEYINPUT113), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n921), .B1(new_n497), .B2(new_n501), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n925), .B1(new_n954), .B2(new_n923), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n840), .A2(new_n957), .A3(KEYINPUT45), .A4(new_n921), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n831), .A2(KEYINPUT45), .A3(new_n839), .A4(new_n921), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(G1971), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n835), .B2(new_n838), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n966), .A3(new_n926), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(G2090), .ZN(new_n968));
  OAI211_X1 g543(.A(G8), .B(new_n953), .C1(new_n962), .C2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(G8), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n964), .B2(new_n926), .ZN(new_n971));
  INV_X1    g546(.A(G1976), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(G288), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n674), .A2(G1976), .ZN(new_n974));
  OR3_X1    g549(.A1(new_n973), .A2(KEYINPUT52), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(KEYINPUT52), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT115), .B(G1981), .Z(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n569), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1981), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n569), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT49), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n971), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n975), .A2(new_n976), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n955), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n681), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n926), .B1(new_n964), .B2(new_n965), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT117), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(new_n926), .C1(new_n964), .C2(new_n965), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(G2090), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n969), .B(new_n984), .C1(new_n996), .C2(new_n953), .ZN(new_n997));
  INV_X1    g572(.A(new_n970), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT45), .B(new_n921), .C1(new_n497), .C2(new_n501), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n926), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n835), .A2(new_n838), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n1002), .B2(new_n921), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n999), .B(new_n762), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2084), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n963), .A2(new_n966), .A3(new_n1005), .A4(new_n926), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1000), .B(new_n926), .C1(KEYINPUT45), .C2(new_n964), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n999), .B1(new_n1008), .B2(new_n762), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G286), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n948), .B1(new_n997), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT120), .B(new_n948), .C1(new_n997), .C2(new_n1011), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT63), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n984), .A2(KEYINPUT116), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n975), .A2(new_n976), .A3(new_n983), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1016), .B(new_n1011), .C1(new_n1017), .C2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n962), .B2(new_n968), .ZN(new_n1022));
  INV_X1    g597(.A(new_n953), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n969), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1014), .A2(new_n1015), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n961), .A2(G1971), .B1(new_n994), .B2(G2090), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n998), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1018), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G2078), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n926), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n922), .B2(new_n923), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT125), .B(new_n1033), .C1(new_n985), .C2(new_n986), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n967), .A2(new_n779), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n958), .A2(new_n960), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT125), .B1(new_n1037), .B2(new_n1033), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1030), .B1(new_n987), .B2(G2078), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n531), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1008), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1042), .A2(new_n1031), .B1(new_n967), .B2(new_n779), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(G301), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT54), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1029), .B(new_n969), .C1(new_n1041), .C2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n582), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1036), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1038), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(G301), .A4(new_n1040), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1048), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n552), .A2(KEYINPUT57), .ZN(new_n1056));
  AOI22_X1  g631(.A1(G299), .A2(KEYINPUT57), .B1(new_n555), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n955), .B(new_n1058), .C1(new_n985), .C2(new_n986), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n994), .A2(new_n750), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n967), .A2(new_n758), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n964), .A2(new_n926), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(G2067), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1065), .A2(new_n592), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1061), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1062), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1061), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT58), .B(G1341), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT121), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n987), .B2(G1996), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n538), .ZN(new_n1077));
  OR2_X1    g652(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1078));
  NAND2_X1  g653(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1069), .A2(new_n1072), .A3(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1076), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n538), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1065), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1065), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1067), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G168), .A2(new_n970), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1007), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1009), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1010), .A2(KEYINPUT123), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT123), .B1(new_n1010), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1093), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1055), .A2(new_n1088), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1105));
  INV_X1    g680(.A(new_n969), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g682(.A(G1976), .B(G288), .C1(new_n982), .C2(new_n971), .ZN(new_n1108));
  INV_X1    g683(.A(new_n979), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n971), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1026), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1095), .A2(new_n1100), .A3(new_n1096), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n1114), .B2(new_n1093), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1096), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1010), .A2(KEYINPUT123), .A3(new_n1094), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1101), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1093), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n997), .A2(new_n1050), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1115), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT126), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1115), .A2(new_n1122), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT127), .B(new_n947), .C1(new_n1113), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1046), .A2(new_n1102), .A3(new_n1054), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1111), .B1(new_n1130), .B2(new_n1088), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(new_n1026), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT127), .B1(new_n1132), .B2(new_n947), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n945), .B1(new_n1129), .B2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g709(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1136));
  AND3_X1   g710(.A1(new_n1136), .A2(new_n849), .A3(new_n911), .ZN(G308));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n911), .A3(new_n849), .ZN(G225));
endmodule


