

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, n1039, G284, G297, G282, G295, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(G543), .B(KEYINPUT0), .Z(n541) );
  NAND2_X2 U552 ( .A1(n738), .A2(n737), .ZN(n751) );
  AND2_X2 U553 ( .A1(n565), .A2(n564), .ZN(G164) );
  XNOR2_X2 U554 ( .A(n534), .B(n533), .ZN(n576) );
  XNOR2_X2 U555 ( .A(n529), .B(n528), .ZN(n617) );
  XNOR2_X2 U556 ( .A(n527), .B(KEYINPUT17), .ZN(n529) );
  AND2_X1 U557 ( .A1(n524), .A2(G2105), .ZN(n613) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n689) );
  AND2_X1 U559 ( .A1(n530), .A2(n520), .ZN(n531) );
  AND2_X2 U560 ( .A1(n522), .A2(G2104), .ZN(n883) );
  INV_X2 U561 ( .A(KEYINPUT66), .ZN(n527) );
  XNOR2_X1 U562 ( .A(n689), .B(KEYINPUT64), .ZN(n786) );
  AND2_X1 U563 ( .A1(n532), .A2(n531), .ZN(G160) );
  XNOR2_X1 U564 ( .A(n720), .B(KEYINPUT103), .ZN(n721) );
  INV_X1 U565 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U566 ( .A1(n569), .A2(G56), .ZN(n570) );
  INV_X1 U567 ( .A(G2104), .ZN(n524) );
  NOR2_X1 U568 ( .A1(n563), .A2(n519), .ZN(n564) );
  XOR2_X1 U569 ( .A(n757), .B(KEYINPUT106), .Z(n518) );
  NAND2_X2 U570 ( .A1(n1039), .A2(G40), .ZN(n785) );
  NAND2_X1 U571 ( .A1(n562), .A2(n561), .ZN(n519) );
  AND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n520) );
  AND2_X1 U573 ( .A1(G43), .A2(n658), .ZN(n521) );
  NOR2_X2 U574 ( .A1(G543), .A2(G651), .ZN(n572) );
  INV_X1 U575 ( .A(KEYINPUT29), .ZN(n720) );
  INV_X1 U576 ( .A(n778), .ZN(n768) );
  NAND2_X1 U577 ( .A1(n769), .A2(n768), .ZN(n770) );
  INV_X1 U578 ( .A(KEYINPUT12), .ZN(n573) );
  XNOR2_X1 U579 ( .A(n573), .B(KEYINPUT75), .ZN(n574) );
  XNOR2_X1 U580 ( .A(n575), .B(n574), .ZN(n578) );
  INV_X1 U581 ( .A(KEYINPUT68), .ZN(n533) );
  INV_X1 U582 ( .A(KEYINPUT1), .ZN(n543) );
  BUF_X1 U583 ( .A(n613), .Z(n888) );
  XNOR2_X1 U584 ( .A(n544), .B(n543), .ZN(n569) );
  NOR2_X2 U585 ( .A1(G651), .A2(n541), .ZN(n658) );
  AND2_X2 U586 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  BUF_X1 U587 ( .A(n569), .Z(n659) );
  AND2_X2 U588 ( .A1(n532), .A2(n531), .ZN(n1039) );
  NAND2_X1 U589 ( .A1(G101), .A2(n883), .ZN(n523) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n523), .Z(n532) );
  NAND2_X1 U591 ( .A1(G125), .A2(n613), .ZN(n526) );
  NAND2_X1 U592 ( .A1(G113), .A2(n889), .ZN(n525) );
  NOR2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  NAND2_X1 U594 ( .A1(G137), .A2(n617), .ZN(n530) );
  INV_X1 U595 ( .A(G651), .ZN(n542) );
  OR2_X2 U596 ( .A1(n542), .A2(n541), .ZN(n534) );
  BUF_X1 U597 ( .A(n576), .Z(n654) );
  NAND2_X1 U598 ( .A1(n654), .A2(G76), .ZN(n538) );
  XOR2_X1 U599 ( .A(KEYINPUT4), .B(KEYINPUT79), .Z(n536) );
  NAND2_X1 U600 ( .A1(G89), .A2(n572), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT80), .ZN(n540) );
  XNOR2_X1 U604 ( .A(KEYINPUT5), .B(n540), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G51), .A2(n658), .ZN(n546) );
  NOR2_X1 U606 ( .A1(G543), .A2(n542), .ZN(n544) );
  NAND2_X1 U607 ( .A1(G63), .A2(n659), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT81), .B(KEYINPUT7), .Z(n550) );
  XNOR2_X1 U612 ( .A(n551), .B(n550), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G90), .A2(n572), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G77), .A2(n654), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT9), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G64), .A2(n659), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n658), .A2(G52), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT70), .B(n557), .Z(n558) );
  NOR2_X1 U622 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U624 ( .A1(n617), .A2(G138), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n613), .A2(G126), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT91), .B(n560), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G102), .A2(n883), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G114), .A2(n889), .ZN(n561) );
  INV_X1 U629 ( .A(G57), .ZN(G237) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  INV_X1 U631 ( .A(G82), .ZN(G220) );
  XOR2_X1 U632 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n567) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G223) );
  XOR2_X1 U635 ( .A(G223), .B(KEYINPUT74), .Z(n839) );
  NAND2_X1 U636 ( .A1(n839), .A2(G567), .ZN(n568) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  XOR2_X1 U638 ( .A(G860), .B(KEYINPUT77), .Z(n605) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NOR2_X1 U640 ( .A1(n571), .A2(n521), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G81), .A2(n572), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(G68), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT13), .ZN(n580) );
  AND2_X2 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X2 U646 ( .A(n582), .B(KEYINPUT76), .ZN(n998) );
  NAND2_X1 U647 ( .A1(n605), .A2(n998), .ZN(G153) );
  XOR2_X1 U648 ( .A(G171), .B(KEYINPUT78), .Z(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G92), .A2(n572), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G79), .A2(n654), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G54), .A2(n658), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G66), .A2(n659), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT15), .B(n589), .ZN(n983) );
  INV_X1 U658 ( .A(G868), .ZN(n672) );
  NAND2_X1 U659 ( .A1(n983), .A2(n672), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G65), .A2(n659), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G91), .A2(n572), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G78), .A2(n654), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G53), .A2(n658), .ZN(n594) );
  XNOR2_X1 U666 ( .A(KEYINPUT71), .B(n594), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT72), .ZN(G299) );
  XOR2_X1 U670 ( .A(KEYINPUT82), .B(G868), .Z(n600) );
  NOR2_X1 U671 ( .A1(G286), .A2(n600), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT83), .B(n601), .Z(n603) );
  NOR2_X1 U673 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(G297) );
  INV_X1 U675 ( .A(G559), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT84), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n983), .A2(n607), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT16), .B(n608), .Z(G148) );
  INV_X1 U680 ( .A(n998), .ZN(n697) );
  NOR2_X1 U681 ( .A1(n697), .A2(G868), .ZN(n611) );
  INV_X1 U682 ( .A(n983), .ZN(n706) );
  NAND2_X1 U683 ( .A1(n706), .A2(G868), .ZN(n609) );
  NOR2_X1 U684 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U686 ( .A(KEYINPUT85), .B(n612), .Z(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n888), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n883), .A2(G99), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n889), .A2(G111), .ZN(n619) );
  BUF_X1 U692 ( .A(n617), .Z(n884) );
  NAND2_X1 U693 ( .A1(G135), .A2(n884), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n939) );
  XNOR2_X1 U696 ( .A(n939), .B(G2096), .ZN(n622) );
  INV_X1 U697 ( .A(G2100), .ZN(n847) );
  NAND2_X1 U698 ( .A1(n622), .A2(n847), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n706), .ZN(n623) );
  XOR2_X1 U700 ( .A(n623), .B(n998), .Z(n669) );
  XNOR2_X1 U701 ( .A(KEYINPUT86), .B(n669), .ZN(n624) );
  NOR2_X1 U702 ( .A1(G860), .A2(n624), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G93), .A2(n572), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G55), .A2(n658), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G80), .A2(n654), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT87), .B(n627), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n659), .A2(G67), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n671) );
  XOR2_X1 U711 ( .A(n632), .B(n671), .Z(G145) );
  NAND2_X1 U712 ( .A1(G49), .A2(n658), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n659), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n541), .A2(G87), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G88), .A2(n572), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G75), .A2(n654), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G50), .A2(n658), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G62), .A2(n659), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G166) );
  INV_X1 U725 ( .A(G166), .ZN(G303) );
  NAND2_X1 U726 ( .A1(G61), .A2(n659), .ZN(n644) );
  XNOR2_X1 U727 ( .A(n644), .B(KEYINPUT88), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G73), .A2(n654), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n645), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G48), .A2(n658), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G86), .A2(n572), .ZN(n648) );
  XNOR2_X1 U733 ( .A(KEYINPUT89), .B(n648), .ZN(n649) );
  NOR2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U736 ( .A1(n572), .A2(G85), .ZN(n653) );
  XOR2_X1 U737 ( .A(KEYINPUT67), .B(n653), .Z(n656) );
  NAND2_X1 U738 ( .A1(G72), .A2(n654), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U740 ( .A(KEYINPUT69), .B(n657), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G47), .A2(n658), .ZN(n661) );
  NAND2_X1 U742 ( .A1(G60), .A2(n659), .ZN(n660) );
  AND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(G290) );
  XNOR2_X1 U745 ( .A(G299), .B(KEYINPUT19), .ZN(n665) );
  XOR2_X1 U746 ( .A(G288), .B(G303), .Z(n664) );
  XNOR2_X1 U747 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(G305), .ZN(n667) );
  XNOR2_X1 U749 ( .A(n667), .B(n671), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(G290), .ZN(n910) );
  XNOR2_X1 U751 ( .A(n910), .B(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT90), .B(n679), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U764 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G96), .A2(n682), .ZN(n844) );
  NAND2_X1 U766 ( .A1(n844), .A2(G2106), .ZN(n686) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U768 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G108), .A2(n684), .ZN(n845) );
  NAND2_X1 U770 ( .A1(n845), .A2(G567), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n846) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n846), .A2(n687), .ZN(n843) );
  NAND2_X1 U774 ( .A1(n843), .A2(G36), .ZN(G176) );
  XNOR2_X1 U775 ( .A(n785), .B(KEYINPUT97), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n786), .A2(n690), .ZN(n693) );
  INV_X1 U777 ( .A(G1996), .ZN(n856) );
  NOR2_X2 U778 ( .A1(n693), .A2(n856), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n691), .B(KEYINPUT26), .ZN(n692) );
  INV_X1 U780 ( .A(n692), .ZN(n695) );
  BUF_X2 U781 ( .A(n693), .Z(n739) );
  NAND2_X1 U782 ( .A1(n739), .A2(G1341), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n699) );
  INV_X1 U785 ( .A(KEYINPUT65), .ZN(n698) );
  XNOR2_X1 U786 ( .A(n699), .B(n698), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n705), .A2(n706), .ZN(n703) );
  INV_X1 U788 ( .A(n739), .ZN(n724) );
  NOR2_X1 U789 ( .A1(n724), .A2(G1348), .ZN(n701) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n739), .ZN(n700) );
  NOR2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(KEYINPUT101), .ZN(n708) );
  NOR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n714) );
  INV_X1 U796 ( .A(G2072), .ZN(n963) );
  NOR2_X1 U797 ( .A1(n739), .A2(n963), .ZN(n710) );
  XNOR2_X1 U798 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n709) );
  XNOR2_X1 U799 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n739), .A2(G1956), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U802 ( .A1(G299), .A2(n716), .ZN(n713) );
  NOR2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U804 ( .A(KEYINPUT102), .B(n715), .ZN(n719) );
  NAND2_X1 U805 ( .A1(G299), .A2(n716), .ZN(n717) );
  XOR2_X1 U806 ( .A(n717), .B(KEYINPUT28), .Z(n718) );
  NOR2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n722) );
  XNOR2_X1 U808 ( .A(n722), .B(n721), .ZN(n729) );
  NOR2_X1 U809 ( .A1(n724), .A2(G1961), .ZN(n723) );
  XOR2_X1 U810 ( .A(KEYINPUT98), .B(n723), .Z(n726) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n959) );
  NAND2_X1 U812 ( .A1(n724), .A2(n959), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n733) );
  NAND2_X1 U814 ( .A1(G171), .A2(n733), .ZN(n727) );
  XOR2_X1 U815 ( .A(KEYINPUT99), .B(n727), .Z(n728) );
  NAND2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n738) );
  NAND2_X1 U817 ( .A1(n739), .A2(G8), .ZN(n778) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n778), .ZN(n753) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n739), .ZN(n749) );
  NOR2_X1 U820 ( .A1(n753), .A2(n749), .ZN(n730) );
  NAND2_X1 U821 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U823 ( .A1(G168), .A2(n732), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G171), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U827 ( .A1(n751), .A2(G286), .ZN(n744) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n778), .ZN(n741) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT104), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n746), .A2(G8), .ZN(n748) );
  INV_X1 U835 ( .A(KEYINPUT32), .ZN(n747) );
  XNOR2_X1 U836 ( .A(n748), .B(n747), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n761) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G8), .A2(n756), .ZN(n757) );
  OR2_X2 U843 ( .A1(n761), .A2(n518), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n758), .A2(n778), .ZN(n760) );
  INV_X1 U845 ( .A(KEYINPUT107), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n760), .B(n759), .ZN(n784) );
  OR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n763) );
  INV_X1 U848 ( .A(G1971), .ZN(n988) );
  NAND2_X1 U849 ( .A1(G166), .A2(n988), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n994) );
  NOR2_X1 U851 ( .A1(n761), .A2(n994), .ZN(n771) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n991) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n773) );
  OR2_X1 U854 ( .A1(n778), .A2(n763), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n773), .A2(n764), .ZN(n765) );
  XNOR2_X1 U856 ( .A(n765), .B(KEYINPUT105), .ZN(n772) );
  AND2_X1 U857 ( .A1(n991), .A2(n772), .ZN(n767) );
  XNOR2_X1 U858 ( .A(G1981), .B(G305), .ZN(n1002) );
  INV_X1 U859 ( .A(n1002), .ZN(n766) );
  AND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n782) );
  INV_X1 U862 ( .A(n772), .ZN(n774) );
  OR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U864 ( .A1(n1002), .A2(n775), .ZN(n780) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U866 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n821) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n834) );
  NAND2_X1 U872 ( .A1(G128), .A2(n888), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G116), .A2(n889), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n789), .B(KEYINPUT35), .ZN(n794) );
  NAND2_X1 U876 ( .A1(G104), .A2(n883), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G140), .A2(n884), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT34), .B(n792), .Z(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U881 ( .A(n795), .B(KEYINPUT36), .Z(n899) );
  XNOR2_X1 U882 ( .A(KEYINPUT37), .B(G2067), .ZN(n831) );
  NOR2_X1 U883 ( .A1(n899), .A2(n831), .ZN(n931) );
  NAND2_X1 U884 ( .A1(n834), .A2(n931), .ZN(n829) );
  INV_X1 U885 ( .A(n829), .ZN(n819) );
  NAND2_X1 U886 ( .A1(G119), .A2(n888), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G131), .A2(n884), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G95), .A2(n883), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G107), .A2(n889), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U893 ( .A(KEYINPUT92), .B(n802), .Z(n906) );
  NAND2_X1 U894 ( .A1(n906), .A2(G1991), .ZN(n813) );
  NAND2_X1 U895 ( .A1(G105), .A2(n883), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT93), .B(n803), .Z(n804) );
  XNOR2_X1 U897 ( .A(n804), .B(KEYINPUT38), .ZN(n806) );
  NAND2_X1 U898 ( .A1(G129), .A2(n888), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n889), .A2(G117), .ZN(n808) );
  NAND2_X1 U901 ( .A1(G141), .A2(n884), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U904 ( .A(KEYINPUT94), .B(n811), .Z(n905) );
  NAND2_X1 U905 ( .A1(n905), .A2(G1996), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT95), .B(n814), .Z(n941) );
  NAND2_X1 U908 ( .A1(n941), .A2(n834), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT96), .ZN(n817) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U911 ( .A1(n987), .A2(n834), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT108), .ZN(n836) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n905), .ZN(n935) );
  NOR2_X1 U917 ( .A1(n906), .A2(G1991), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT110), .ZN(n940) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n824) );
  XOR2_X1 U920 ( .A(n824), .B(KEYINPUT109), .Z(n825) );
  NOR2_X1 U921 ( .A1(n940), .A2(n825), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n826), .A2(n941), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n935), .A2(n827), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(KEYINPUT39), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n899), .A2(n831), .ZN(n933) );
  NAND2_X1 U927 ( .A1(n832), .A2(n933), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n838) );
  XOR2_X1 U930 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n837) );
  XNOR2_X1 U931 ( .A(n838), .B(n837), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  XOR2_X1 U936 ( .A(KEYINPUT113), .B(n841), .Z(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  INV_X1 U944 ( .A(n846), .ZN(G319) );
  XNOR2_X1 U945 ( .A(n847), .B(G2096), .ZN(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XOR2_X1 U949 ( .A(G2067), .B(n963), .Z(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U954 ( .A(KEYINPUT41), .B(G1961), .Z(n858) );
  XOR2_X1 U955 ( .A(n856), .B(G1991), .Z(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n859), .B(KEYINPUT115), .Z(n861) );
  XOR2_X1 U958 ( .A(G1976), .B(n988), .Z(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U960 ( .A(G1956), .B(G1966), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1981), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT114), .B(G2474), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n888), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n883), .A2(G100), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n889), .A2(G112), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G136), .A2(n884), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G103), .A2(n883), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G139), .A2(n884), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G127), .A2(n888), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G115), .A2(n889), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(KEYINPUT117), .B(n879), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT47), .B(n880), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n944) );
  NAND2_X1 U983 ( .A1(G106), .A2(n883), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G142), .A2(n884), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(KEYINPUT45), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(KEYINPUT116), .B(n892), .Z(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n895), .B(G162), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n944), .B(n896), .ZN(n904) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  XNOR2_X1 U995 ( .A(n939), .B(KEYINPUT118), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U998 ( .A(G160), .B(G164), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1004 ( .A(n910), .B(G286), .Z(n912) );
  XOR2_X1 U1005 ( .A(n983), .B(G171), .Z(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1007 ( .A(n913), .B(n998), .Z(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G397) );
  XOR2_X1 U1009 ( .A(G2438), .B(G2435), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2430), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n917), .B(G2454), .Z(n919) );
  XNOR2_X1 U1013 ( .A(G1341), .B(G1348), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n923) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2427), .Z(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT112), .B(G2446), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1018 ( .A(n923), .B(n922), .Z(n924) );
  NAND2_X1 U1019 ( .A1(G14), .A2(n924), .ZN(n930) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  INV_X1 U1028 ( .A(n930), .ZN(G401) );
  INV_X1 U1029 ( .A(n931), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n954) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n936), .Z(n952) );
  XNOR2_X1 U1034 ( .A(G160), .B(G2084), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n937), .B(KEYINPUT119), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n946) );
  XOR2_X1 U1040 ( .A(G2072), .B(n944), .Z(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT50), .B(n947), .Z(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n948), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n978), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G29), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT121), .B(n958), .Z(n1036) );
  XOR2_X1 U1052 ( .A(n959), .B(G27), .Z(n961) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n965) );
  XOR2_X1 U1058 ( .A(n963), .B(G33), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT122), .B(n966), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT53), .ZN(n974) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G35), .B(G2090), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n978), .B(n977), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(G29), .A2(n979), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n980), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(G11), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n982), .B(KEYINPUT124), .ZN(n1034) );
  INV_X1 U1074 ( .A(G16), .ZN(n1030) );
  XOR2_X1 U1075 ( .A(n1030), .B(KEYINPUT56), .Z(n1008) );
  XNOR2_X1 U1076 ( .A(G171), .B(G1961), .ZN(n985) );
  XOR2_X1 U1077 ( .A(n983), .B(G1348), .Z(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n997) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G299), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n988), .A2(G166), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(KEYINPUT125), .B(n995), .Z(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(n998), .B(G1341), .Z(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(G1966), .B(G168), .Z(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT57), .B(n1003), .Z(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1006), .B(KEYINPUT126), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1032) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1010) );
  XOR2_X1 U1096 ( .A(G1971), .B(G22), .Z(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G24), .B(G1986), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1961), .B(G5), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1027) );
  XOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G4), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G20), .B(G1956), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(G1981), .B(G6), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G1341), .B(G19), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT60), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1119 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1120 ( .A(n1037), .B(KEYINPUT127), .ZN(n1038) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1038), .Z(G150) );
  INV_X1 U1122 ( .A(G150), .ZN(G311) );
endmodule

