

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XOR2_X1 U325 ( .A(n424), .B(n352), .Z(n293) );
  XOR2_X1 U326 ( .A(KEYINPUT25), .B(n409), .Z(n294) );
  XNOR2_X1 U327 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n455) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U329 ( .A(KEYINPUT96), .ZN(n412) );
  XNOR2_X1 U330 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U331 ( .A(G57GAT), .B(KEYINPUT13), .Z(n439) );
  XNOR2_X1 U332 ( .A(n442), .B(n441), .ZN(n443) );
  NOR2_X1 U333 ( .A1(n584), .A2(n482), .ZN(n417) );
  NAND2_X1 U334 ( .A1(n414), .A2(n534), .ZN(n415) );
  XNOR2_X1 U335 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U336 ( .A(KEYINPUT94), .ZN(n355) );
  XNOR2_X1 U337 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U338 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U339 ( .A1(n476), .A2(n475), .ZN(n570) );
  INV_X1 U340 ( .A(G99GAT), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n364), .B(n381), .ZN(n523) );
  XNOR2_X1 U342 ( .A(n477), .B(G176GAT), .ZN(n478) );
  XNOR2_X1 U343 ( .A(n452), .B(KEYINPUT112), .ZN(n453) );
  XNOR2_X1 U344 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n454), .B(n453), .ZN(G1338GAT) );
  XOR2_X1 U346 ( .A(G190GAT), .B(G134GAT), .Z(n323) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n295), .B(G120GAT), .ZN(n438) );
  XOR2_X1 U349 ( .A(n323), .B(n438), .Z(n297) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U352 ( .A(G176GAT), .B(KEYINPUT84), .Z(n299) );
  XNOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U355 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n302), .B(G113GAT), .ZN(n429) );
  XNOR2_X1 U358 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n303), .B(KEYINPUT81), .ZN(n395) );
  XNOR2_X1 U360 ( .A(n429), .B(n395), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT17), .B(G183GAT), .Z(n307) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U365 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n308) );
  XOR2_X1 U366 ( .A(n309), .B(n308), .Z(n360) );
  XNOR2_X1 U367 ( .A(n310), .B(n360), .ZN(n535) );
  INV_X1 U368 ( .A(n535), .ZN(n476) );
  XOR2_X1 U369 ( .A(KEYINPUT7), .B(G50GAT), .Z(n312) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(G29GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U372 ( .A(KEYINPUT8), .B(n313), .Z(n423) );
  XOR2_X1 U373 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n315) );
  XNOR2_X1 U374 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n423), .B(n316), .ZN(n327) );
  XOR2_X1 U377 ( .A(G85GAT), .B(G92GAT), .Z(n442) );
  XOR2_X1 U378 ( .A(KEYINPUT72), .B(G162GAT), .Z(n367) );
  XOR2_X1 U379 ( .A(n442), .B(n367), .Z(n318) );
  XNOR2_X1 U380 ( .A(G218GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U382 ( .A(KEYINPUT74), .B(G99GAT), .Z(n320) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U385 ( .A(n322), .B(n321), .Z(n325) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n569) );
  XNOR2_X1 U389 ( .A(n569), .B(KEYINPUT101), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n328), .B(KEYINPUT36), .ZN(n587) );
  XOR2_X1 U391 ( .A(KEYINPUT76), .B(KEYINPUT80), .Z(n330) );
  XNOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n349) );
  XOR2_X1 U394 ( .A(G71GAT), .B(G127GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U397 ( .A(KEYINPUT75), .B(G64GAT), .Z(n334) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G1GAT), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U400 ( .A(n336), .B(n335), .Z(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n338) );
  XNOR2_X1 U402 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n345) );
  XOR2_X1 U404 ( .A(G155GAT), .B(G78GAT), .Z(n340) );
  XNOR2_X1 U405 ( .A(G22GAT), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U407 ( .A(n439), .B(n341), .Z(n343) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n349), .B(n348), .Z(n559) );
  INV_X1 U413 ( .A(n559), .ZN(n584) );
  XOR2_X1 U414 ( .A(G197GAT), .B(G8GAT), .Z(n424) );
  XOR2_X1 U415 ( .A(KEYINPUT93), .B(G92GAT), .Z(n351) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  NAND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n293), .B(n353), .ZN(n358) );
  XNOR2_X1 U420 ( .A(G176GAT), .B(G204GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n354), .B(G64GAT), .ZN(n437) );
  XNOR2_X1 U422 ( .A(n437), .B(KEYINPUT95), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT21), .B(G218GAT), .Z(n362) );
  XNOR2_X1 U425 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(KEYINPUT87), .B(n363), .ZN(n381) );
  XNOR2_X1 U428 ( .A(KEYINPUT27), .B(n523), .ZN(n531) );
  XOR2_X1 U429 ( .A(G155GAT), .B(KEYINPUT2), .Z(n366) );
  XNOR2_X1 U430 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n402) );
  XOR2_X1 U432 ( .A(n402), .B(n367), .Z(n373) );
  XOR2_X1 U433 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U434 ( .A(G106GAT), .B(G78GAT), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n368), .B(G148GAT), .ZN(n446) );
  XOR2_X1 U436 ( .A(KEYINPUT86), .B(n446), .Z(n370) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n425), .B(n371), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n375) );
  XNOR2_X1 U442 ( .A(G50GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U444 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n379) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(KEYINPUT24), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U448 ( .A(n381), .B(n380), .Z(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n472) );
  XOR2_X1 U450 ( .A(n472), .B(KEYINPUT64), .Z(n384) );
  XNOR2_X1 U451 ( .A(KEYINPUT28), .B(n384), .ZN(n537) );
  XNOR2_X1 U452 ( .A(KEYINPUT85), .B(n476), .ZN(n385) );
  NOR2_X1 U453 ( .A1(n537), .A2(n385), .ZN(n386) );
  NAND2_X1 U454 ( .A1(n531), .A2(n386), .ZN(n407) );
  XOR2_X1 U455 ( .A(KEYINPUT6), .B(G57GAT), .Z(n388) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n388), .B(n387), .ZN(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT74), .B(G162GAT), .Z(n390) );
  XNOR2_X1 U459 ( .A(G141GAT), .B(G134GAT), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(G148GAT), .Z(n392) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U463 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U464 ( .A(n394), .B(n393), .Z(n400) );
  XOR2_X1 U465 ( .A(G85GAT), .B(n395), .Z(n397) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(n398), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U470 ( .A(n401), .B(KEYINPUT4), .Z(n404) );
  XNOR2_X1 U471 ( .A(n402), .B(KEYINPUT5), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U473 ( .A(n406), .B(n405), .Z(n510) );
  NAND2_X1 U474 ( .A1(n407), .A2(n510), .ZN(n416) );
  NAND2_X1 U475 ( .A1(n535), .A2(n523), .ZN(n408) );
  NAND2_X1 U476 ( .A1(n472), .A2(n408), .ZN(n409) );
  NOR2_X1 U477 ( .A1(n472), .A2(n535), .ZN(n410) );
  XNOR2_X1 U478 ( .A(KEYINPUT26), .B(n410), .ZN(n574) );
  NAND2_X1 U479 ( .A1(n531), .A2(n574), .ZN(n411) );
  NAND2_X1 U480 ( .A1(n294), .A2(n411), .ZN(n413) );
  INV_X1 U481 ( .A(n510), .ZN(n534) );
  NAND2_X1 U482 ( .A1(n416), .A2(n415), .ZN(n482) );
  XOR2_X1 U483 ( .A(KEYINPUT102), .B(n417), .Z(n418) );
  NOR2_X1 U484 ( .A1(n587), .A2(n418), .ZN(n419) );
  XNOR2_X1 U485 ( .A(KEYINPUT37), .B(n419), .ZN(n495) );
  XOR2_X1 U486 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n421) );
  XNOR2_X1 U487 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT65), .B(KEYINPUT69), .Z(n427) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n428), .B(G1GAT), .Z(n434) );
  XOR2_X1 U494 ( .A(n429), .B(KEYINPUT29), .Z(n431) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n576) );
  INV_X1 U500 ( .A(n576), .ZN(n551) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n439), .B(KEYINPUT31), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n440), .B(KEYINPUT33), .ZN(n444) );
  AND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XOR2_X1 U505 ( .A(KEYINPUT32), .B(n445), .Z(n448) );
  XNOR2_X1 U506 ( .A(n446), .B(KEYINPUT71), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n461) );
  XOR2_X1 U509 ( .A(n461), .B(KEYINPUT41), .Z(n556) );
  INV_X1 U510 ( .A(n556), .ZN(n540) );
  NAND2_X1 U511 ( .A1(n551), .A2(n540), .ZN(n508) );
  NOR2_X1 U512 ( .A1(n495), .A2(n508), .ZN(n451) );
  XOR2_X1 U513 ( .A(KEYINPUT110), .B(n451), .Z(n526) );
  NOR2_X1 U514 ( .A1(n476), .A2(n526), .ZN(n454) );
  INV_X1 U515 ( .A(n569), .ZN(n563) );
  OR2_X1 U516 ( .A1(n556), .A2(n551), .ZN(n456) );
  AND2_X1 U517 ( .A1(n457), .A2(n559), .ZN(n458) );
  AND2_X1 U518 ( .A1(n563), .A2(n458), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT47), .B(n459), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n587), .A2(n559), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT45), .B(n460), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT115), .B(n463), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT70), .B(n551), .Z(n566) );
  INV_X1 U525 ( .A(n566), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT48), .ZN(n532) );
  NAND2_X1 U529 ( .A1(n532), .A2(n523), .ZN(n470) );
  XOR2_X1 U530 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n510), .A2(n471), .ZN(n573) );
  NAND2_X1 U533 ( .A1(n573), .A2(n472), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT124), .B(KEYINPUT55), .Z(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n570), .A2(n540), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n477) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  NOR2_X1 U539 ( .A1(n569), .A2(n559), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT97), .B(n483), .ZN(n507) );
  NAND2_X1 U543 ( .A1(n461), .A2(n566), .ZN(n494) );
  NOR2_X1 U544 ( .A1(n507), .A2(n494), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT98), .ZN(n491) );
  NAND2_X1 U546 ( .A1(n510), .A2(n491), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n491), .A2(n523), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U551 ( .A1(n491), .A2(n535), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NAND2_X1 U554 ( .A1(n491), .A2(n537), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT100), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NOR2_X1 U558 ( .A1(n495), .A2(n494), .ZN(n497) );
  XOR2_X1 U559 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n505) );
  NAND2_X1 U561 ( .A1(n510), .A2(n505), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n505), .A2(n523), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U567 ( .A1(n505), .A2(n535), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n505), .A2(n537), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n512) );
  NOR2_X1 U573 ( .A1(n508), .A2(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(KEYINPUT107), .B(n509), .Z(n518) );
  NAND2_X1 U575 ( .A1(n518), .A2(n510), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NAND2_X1 U578 ( .A1(n523), .A2(n518), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U581 ( .A1(n518), .A2(n535), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n537), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n526), .A2(n534), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  INV_X1 U590 ( .A(n523), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n524), .A2(n526), .ZN(n525) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n529) );
  INV_X1 U594 ( .A(n537), .ZN(n527) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n550), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT116), .B(n536), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n566), .A2(n545), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n584), .A2(n545), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n569), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT118), .Z(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n574), .ZN(n562) );
  NOR2_X1 U617 ( .A1(n551), .A2(n562), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n556), .A2(n562), .ZN(n557) );
  XOR2_X1 U624 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n562), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n564), .Z(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT122), .B(n565), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n570), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n584), .A2(n570), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G190GAT), .ZN(G1351GAT) );
  AND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT125), .ZN(n586) );
  INV_X1 U640 ( .A(n586), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n583), .A2(n576), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  OR2_X1 U647 ( .A1(n586), .A2(n461), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

