//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  NOR2_X1   g0019(.A1(new_n206), .A2(new_n207), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n211), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n219), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  INV_X1    g0037(.A(G107), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G97), .ZN(new_n239));
  INV_X1    g0039(.A(G97), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G107), .ZN(new_n241));
  AND2_X1   g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n207), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G33), .A3(G41), .ZN(new_n258));
  INV_X1    g0058(.A(new_n221), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(new_n252), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT67), .A3(G222), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n264), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n273), .A2(G223), .B1(G77), .B2(new_n272), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  INV_X1    g0075(.A(G222), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n267), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n254), .B(new_n262), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .A3(new_n221), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT68), .B1(new_n283), .B2(new_n221), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT8), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n288), .A2(KEYINPUT69), .A3(G58), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(G58), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT69), .B1(new_n288), .B2(G58), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n222), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n222), .A2(new_n268), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n292), .A2(new_n294), .B1(G150), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n208), .A2(G20), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n287), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n286), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n284), .C1(G1), .C2(new_n222), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(new_n207), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n282), .B1(G169), .B2(new_n280), .C1(new_n299), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n299), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT71), .ZN(new_n308));
  INV_X1    g0108(.A(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT71), .B1(new_n299), .B2(new_n305), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT72), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n280), .A2(G190), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n280), .A2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n314), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n306), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n254), .B1(new_n261), .B2(G232), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n263), .A2(G226), .A3(G1698), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n269), .A2(new_n271), .A3(G223), .A4(new_n264), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G87), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n279), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n324), .A2(G179), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n324), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G159), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n295), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G58), .A2(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n203), .A2(new_n205), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(new_n337), .B2(G20), .ZN(new_n338));
  AOI21_X1  g0138(.A(G20), .B1(new_n269), .B2(new_n271), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n272), .A2(new_n342), .A3(new_n222), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT16), .B(new_n338), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n342), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(G68), .C1(new_n340), .C2(new_n339), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT16), .A4(new_n338), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n272), .A2(new_n222), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n340), .B(G20), .C1(new_n269), .C2(new_n271), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n338), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n287), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n304), .A2(new_n292), .ZN(new_n360));
  INV_X1    g0160(.A(new_n300), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n292), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n333), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT18), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  INV_X1    g0166(.A(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n350), .B2(new_n358), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(new_n333), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n324), .A2(G190), .A3(new_n329), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n318), .B1(new_n324), .B2(new_n329), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n359), .A2(new_n373), .A3(new_n363), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT17), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n368), .A2(new_n376), .A3(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n303), .A2(new_n284), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n202), .A2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(G77), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n382), .B1(new_n293), .B2(new_n383), .C1(new_n207), .C2(new_n295), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT75), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n300), .A2(G68), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT12), .ZN(new_n390));
  INV_X1    g0190(.A(new_n304), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n386), .B2(new_n387), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n269), .A2(new_n271), .A3(G226), .A4(new_n264), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT73), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n395), .A2(KEYINPUT73), .A3(new_n396), .A4(new_n397), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n279), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n254), .B1(new_n261), .B2(G238), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n402), .A2(new_n405), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  OAI211_X1 g0208(.A(G190), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n404), .B1(new_n402), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n394), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n410), .B2(new_n411), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(G169), .C1(new_n410), .C2(new_n411), .ZN(new_n417));
  OAI211_X1 g0217(.A(G179), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n394), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n261), .A2(G244), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n266), .A2(KEYINPUT70), .A3(G232), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n273), .A2(G238), .B1(G107), .B2(new_n272), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  INV_X1    g0225(.A(G232), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n265), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n254), .B(new_n422), .C1(new_n428), .C2(new_n279), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n429), .A2(new_n281), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G20), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT8), .B(G58), .ZN(new_n432));
  OR2_X1    g0232(.A1(KEYINPUT15), .A2(G87), .ZN(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT15), .A2(G87), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n431), .B1(new_n432), .B2(new_n295), .C1(new_n293), .C2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n381), .B1(new_n383), .B2(new_n361), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n383), .B2(new_n304), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n429), .B2(G169), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n429), .B2(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n318), .B2(new_n429), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n380), .A2(new_n421), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n323), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT6), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n239), .A2(new_n241), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n238), .A2(KEYINPUT6), .A3(G97), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n450), .A2(new_n222), .B1(new_n383), .B2(new_n295), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n342), .B1(new_n263), .B2(G20), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n238), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n381), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n251), .A2(G33), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n300), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(new_n303), .A3(G97), .A4(new_n284), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G97), .B2(new_n300), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n264), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n279), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n221), .B1(KEYINPUT66), .B2(new_n255), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n258), .A2(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n251), .A2(G45), .A3(G274), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT80), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n477), .A2(G257), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n472), .A2(G179), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n331), .B1(new_n472), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n462), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT82), .B(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n300), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n285), .A2(new_n457), .A3(new_n286), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n283), .A2(new_n221), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n492), .B2(new_n222), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n222), .B1(new_n240), .B2(G33), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n464), .B2(new_n465), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(G20), .B1(new_n221), .B2(new_n283), .ZN(new_n506));
  INV_X1    g0306(.A(new_n498), .ZN(new_n507));
  INV_X1    g0307(.A(new_n465), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n463), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT20), .ZN(new_n510));
  AOI221_X4 g0310(.A(new_n493), .B1(new_n494), .B2(G116), .C1(new_n500), .C2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n264), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(G303), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n263), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n279), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n484), .A2(new_n487), .ZN(new_n517));
  INV_X1    g0317(.A(new_n476), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n260), .B(G270), .C1(new_n482), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(G190), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n511), .B(new_n521), .C1(new_n522), .C2(new_n520), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n353), .B2(new_n354), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n448), .A2(new_n449), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n460), .B1(new_n527), .B2(new_n381), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n472), .A2(G190), .A3(new_n488), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n318), .B1(new_n472), .B2(new_n488), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT81), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n491), .B(new_n523), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n264), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(G1698), .ZN(new_n537));
  INV_X1    g0337(.A(G294), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n268), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n279), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n477), .A2(G264), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n517), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT87), .B1(new_n542), .B2(G190), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n318), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n539), .A2(new_n279), .B1(new_n477), .B2(G264), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n522), .A4(new_n517), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n300), .A2(G107), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT25), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n287), .A2(new_n458), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n238), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n238), .A2(G20), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT23), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT86), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n502), .A2(new_n504), .A3(G33), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(G20), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n222), .A4(G33), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n269), .A2(new_n271), .A3(new_n222), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n263), .A2(new_n562), .A3(new_n222), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n287), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(KEYINPUT24), .A3(new_n564), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n552), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n548), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n535), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n500), .A2(new_n510), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n494), .A2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(new_n493), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n520), .A3(G169), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n516), .A2(G179), .A3(new_n517), .A4(new_n519), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n511), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n575), .A2(new_n520), .A3(KEYINPUT21), .A4(G169), .ZN(new_n582));
  INV_X1    g0382(.A(new_n580), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n575), .A3(KEYINPUT85), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n578), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n542), .A2(new_n331), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G179), .B2(new_n542), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n569), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n476), .B1(new_n473), .B2(new_n258), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n485), .B1(new_n590), .B2(G250), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n269), .A2(new_n271), .A3(G238), .A4(new_n264), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(G1698), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n556), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n279), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n591), .A2(new_n595), .A3(G190), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n318), .B1(new_n591), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n222), .B1(new_n396), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n240), .A3(new_n238), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n269), .A2(new_n271), .A3(new_n222), .A4(G68), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n599), .B1(new_n293), .B2(new_n240), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n381), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n300), .B1(new_n433), .B2(new_n434), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT83), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n607), .A2(new_n612), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n494), .A2(G87), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n598), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n591), .A2(new_n595), .A3(new_n281), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(G169), .B1(new_n591), .B2(new_n595), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n551), .A2(new_n435), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n612), .B1(new_n607), .B2(new_n609), .ZN(new_n623));
  AOI211_X1 g0423(.A(KEYINPUT83), .B(new_n608), .C1(new_n606), .C2(new_n381), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n616), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n616), .B2(new_n626), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n446), .A2(new_n571), .A3(new_n589), .A4(new_n630), .ZN(G372));
  OR2_X1    g0431(.A1(new_n321), .A2(new_n322), .ZN(new_n632));
  INV_X1    g0432(.A(new_n370), .ZN(new_n633));
  INV_X1    g0433(.A(new_n413), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n440), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n419), .A2(new_n420), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n375), .B2(new_n377), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n632), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n306), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n260), .B(G257), .C1(new_n482), .C2(new_n518), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n517), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n468), .A2(new_n469), .ZN(new_n642));
  INV_X1    g0442(.A(new_n469), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n263), .A2(G244), .A3(new_n264), .A4(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n644), .A3(new_n466), .A4(new_n467), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n279), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT81), .B1(new_n646), .B2(new_n318), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(new_n528), .A3(new_n533), .A4(new_n529), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n491), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n611), .A2(new_n613), .B1(G87), .B2(new_n494), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n650), .A2(new_n598), .B1(new_n620), .B2(new_n625), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n548), .A2(new_n569), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n589), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n621), .B1(new_n611), .B2(new_n613), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n594), .A2(new_n279), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n260), .A2(G250), .A3(new_n518), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n483), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n331), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n617), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n615), .B1(new_n623), .B2(new_n624), .ZN(new_n661));
  OAI21_X1  g0461(.A(G200), .B1(new_n656), .B2(new_n658), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n591), .A2(new_n595), .A3(G190), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n655), .A2(new_n660), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT84), .ZN(new_n666));
  INV_X1    g0466(.A(new_n491), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n616), .A2(new_n626), .A3(new_n627), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(new_n626), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT88), .B1(new_n489), .B2(new_n490), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n472), .A2(G179), .A3(new_n488), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n673), .B(new_n674), .C1(new_n646), .C2(new_n331), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n675), .A3(new_n462), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n665), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n654), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n674), .B1(new_n646), .B2(new_n331), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n528), .B1(new_n683), .B2(KEYINPUT88), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n651), .A2(new_n684), .A3(new_n678), .A4(new_n675), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n626), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(KEYINPUT26), .B2(new_n669), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n446), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n639), .A2(new_n690), .ZN(G369));
  AND2_X1   g0491(.A1(new_n222), .A2(G13), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n251), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n575), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n585), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n585), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n523), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n698), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n569), .A2(new_n705), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n570), .A2(new_n706), .B1(new_n569), .B2(new_n587), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n588), .A2(new_n705), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n585), .A2(new_n705), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n710), .A2(new_n707), .B1(new_n588), .B2(new_n705), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n225), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n602), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n220), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n718), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n698), .B1(new_n682), .B2(new_n688), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n726));
  NAND2_X1  g0526(.A1(new_n669), .A2(new_n678), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n677), .A2(KEYINPUT92), .A3(KEYINPUT26), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n651), .A2(new_n684), .A3(new_n675), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n678), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n589), .A2(new_n649), .ZN(new_n733));
  INV_X1    g0533(.A(new_n653), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n626), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(new_n705), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n725), .A2(new_n726), .B1(new_n737), .B2(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n472), .A2(new_n488), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n591), .B2(new_n595), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n542), .A4(new_n520), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n540), .A2(new_n591), .A3(new_n595), .A4(new_n541), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n739), .A2(new_n742), .A3(new_n580), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n656), .A2(new_n658), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n646), .A2(new_n545), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n746), .A2(new_n747), .A3(new_n580), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT90), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n746), .B2(new_n580), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT90), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n741), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n749), .A2(new_n698), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n630), .A2(new_n571), .A3(new_n589), .A4(new_n705), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(KEYINPUT31), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT31), .B(new_n698), .C1(new_n744), .C2(new_n748), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(G330), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n738), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n723), .B1(new_n761), .B2(G1), .ZN(G364));
  AOI21_X1  g0562(.A(new_n251), .B1(new_n692), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n717), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n704), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n702), .A2(new_n703), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n702), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n259), .B1(new_n222), .B2(G169), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n222), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n318), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n263), .B1(new_n781), .B2(G283), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G329), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n281), .A2(new_n318), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(new_n778), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI211_X1 g0590(.A(new_n782), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n222), .A2(new_n522), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n281), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n778), .A2(new_n793), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G322), .A2(new_n795), .B1(new_n797), .B2(G311), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n792), .A2(new_n779), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n792), .A2(new_n787), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n798), .B1(new_n514), .B2(new_n799), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n222), .B1(new_n783), .B2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n791), .B(new_n803), .C1(G294), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n799), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G87), .A2(new_n807), .B1(new_n788), .B2(G68), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(new_n263), .C1(new_n207), .C2(new_n802), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G58), .A2(new_n795), .B1(new_n781), .B2(G107), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n383), .B2(new_n796), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n784), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n784), .B2(new_n334), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n240), .C2(new_n804), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n809), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n777), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n777), .A2(new_n772), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n263), .A2(G355), .A3(new_n225), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n249), .A2(new_n475), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n716), .A2(new_n263), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n721), .B2(G45), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n819), .B1(G116), .B2(new_n225), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n816), .A2(new_n765), .A3(new_n824), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n767), .A2(new_n769), .B1(new_n773), .B2(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n438), .A2(new_n698), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n443), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n441), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n440), .A2(new_n705), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n724), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n698), .B(new_n831), .C1(new_n682), .C2(new_n688), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n760), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n760), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n837), .A2(new_n766), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n777), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n771), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n765), .B1(new_n842), .B2(G77), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n796), .A2(new_n334), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n789), .A2(new_n845), .B1(new_n846), .B2(new_n794), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(G137), .C2(new_n801), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n263), .B1(new_n799), .B2(new_n207), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n780), .A2(new_n202), .B1(new_n784), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(G58), .C2(new_n805), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G311), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n780), .A2(new_n601), .B1(new_n784), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G283), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n789), .A2(new_n858), .B1(new_n796), .B2(new_n505), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT95), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n802), .A2(new_n514), .B1(new_n799), .B2(new_n238), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n272), .B1(new_n804), .B2(new_n240), .C1(new_n538), .C2(new_n794), .ZN(new_n862));
  OR4_X1    g0662(.A1(new_n857), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n843), .B1(new_n864), .B2(new_n777), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n832), .B2(new_n771), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n840), .A2(new_n866), .ZN(G384));
  XNOR2_X1  g0667(.A(new_n450), .B(KEYINPUT97), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT35), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(G116), .A4(new_n223), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  NAND3_X1  g0673(.A1(new_n220), .A2(G77), .A3(new_n336), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n251), .B(G13), .C1(new_n874), .C2(new_n245), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n338), .B1(new_n341), .B2(new_n343), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n877), .B2(KEYINPUT98), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT98), .B2(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n381), .A3(new_n350), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n363), .ZN(new_n881));
  INV_X1    g0681(.A(new_n696), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n379), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  INV_X1    g0686(.A(new_n333), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n202), .B1(new_n452), .B2(new_n453), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n337), .A2(G20), .ZN(new_n889));
  INV_X1    g0689(.A(new_n335), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n357), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n381), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n349), .B2(new_n345), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n887), .B1(new_n894), .B2(new_n367), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n696), .B(KEYINPUT99), .Z(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n894), .B2(new_n367), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(new_n898), .A3(new_n374), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n881), .B1(new_n887), .B2(new_n882), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n359), .A2(new_n363), .A3(new_n373), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n886), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n886), .A2(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n886), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n900), .A2(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n883), .B1(new_n370), .B2(new_n378), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n420), .A2(new_n698), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n636), .A2(new_n634), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n419), .A2(new_n420), .A3(new_n698), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND4_X1   g0718(.A1(KEYINPUT31), .A2(new_n749), .A3(new_n698), .A4(new_n753), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n832), .B(new_n918), .C1(new_n756), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n368), .A2(new_n376), .A3(new_n373), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n376), .B1(new_n368), .B2(new_n373), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT101), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT101), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n375), .A2(new_n926), .A3(new_n377), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n370), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n898), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n901), .A2(new_n364), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT100), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n368), .B2(new_n896), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n931), .A2(new_n898), .B1(KEYINPUT37), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n899), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n904), .B1(new_n938), .B2(KEYINPUT102), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n931), .A2(KEYINPUT100), .A3(KEYINPUT37), .A4(new_n898), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n899), .A2(new_n935), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n929), .B2(new_n928), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT102), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT38), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n922), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n921), .B1(new_n946), .B2(KEYINPUT40), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT105), .ZN(new_n948));
  INV_X1    g0748(.A(new_n919), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n755), .A2(KEYINPUT31), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n754), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(new_n446), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n703), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n948), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n904), .A2(new_n910), .ZN(new_n955));
  INV_X1    g0755(.A(new_n830), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n918), .C1(new_n834), .C2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n370), .A2(new_n897), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n636), .A2(new_n698), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n944), .B1(new_n943), .B2(KEYINPUT38), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n938), .A2(KEYINPUT102), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT39), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n904), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n955), .A2(KEYINPUT39), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT103), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n967), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n961), .ZN(new_n971));
  INV_X1    g0771(.A(new_n918), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n735), .B1(new_n687), .B2(KEYINPUT89), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n680), .A2(new_n681), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n705), .B(new_n832), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n972), .B1(new_n975), .B2(new_n830), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n958), .B1(new_n976), .B2(new_n955), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT103), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n969), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n954), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n982));
  INV_X1    g0782(.A(new_n726), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n446), .C1(new_n724), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n639), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n251), .B2(new_n692), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n981), .A2(new_n986), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n876), .B1(new_n988), .B2(new_n989), .ZN(G367));
  OAI21_X1  g0790(.A(new_n651), .B1(new_n650), .B2(new_n705), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n671), .A2(new_n661), .A3(new_n698), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n772), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n817), .B1(new_n225), .B2(new_n435), .ZN(new_n996));
  INV_X1    g0796(.A(new_n821), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n236), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n765), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT108), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n802), .A2(new_n856), .B1(new_n780), .B2(new_n240), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G294), .B2(new_n788), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n796), .A2(new_n858), .B1(new_n784), .B2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n263), .B(new_n1004), .C1(G303), .C2(new_n795), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n805), .A2(G107), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT46), .B1(new_n799), .B2(new_n501), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n505), .A2(KEYINPUT46), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n799), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G137), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n794), .A2(new_n845), .B1(new_n784), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n263), .B1(new_n802), .B2(new_n846), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n799), .A2(new_n201), .B1(new_n780), .B2(new_n383), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n804), .A2(new_n202), .ZN(new_n1015));
  OR4_X1    g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n797), .A2(G50), .B1(new_n788), .B2(G159), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT47), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n841), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n995), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n982), .B1(new_n724), .B2(new_n983), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n648), .B(new_n491), .C1(new_n528), .C2(new_n705), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n684), .A2(new_n675), .A3(new_n698), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1026), .B1(new_n714), .B2(new_n1029), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n714), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n714), .A2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1030), .A2(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT107), .B1(new_n1036), .B2(new_n713), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n710), .A2(new_n707), .A3(new_n708), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n704), .A2(new_n711), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n713), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1025), .A2(new_n1037), .A3(new_n759), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1031), .A2(new_n1030), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n712), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(new_n713), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT107), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n761), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n717), .B(KEYINPUT41), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n764), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1029), .B(KEYINPUT106), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n588), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n698), .B1(new_n1052), .B2(new_n491), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n709), .A2(new_n733), .A3(new_n710), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT42), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT43), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n1057), .A3(new_n994), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n994), .A2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1051), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n713), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1062), .B(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1024), .B1(new_n1050), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT110), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT110), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n1024), .C1(new_n1050), .C2(new_n1066), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(G387));
  NAND3_X1  g0871(.A1(new_n713), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n738), .B2(new_n760), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1025), .A2(new_n759), .A3(new_n1040), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n717), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n432), .A2(G50), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n475), .B1(new_n202), .B2(new_n383), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT111), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n719), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(new_n1079), .C2(new_n719), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n821), .C1(new_n233), .C2(new_n475), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n263), .A2(new_n225), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1082), .B1(G107), .B2(new_n225), .C1(new_n719), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n766), .B1(new_n1084), .B2(new_n818), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n772), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n804), .A2(new_n435), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n799), .A2(new_n383), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n263), .B1(new_n780), .B2(new_n240), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G68), .C2(new_n797), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n292), .A2(new_n788), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n794), .A2(new_n207), .B1(new_n784), .B2(new_n845), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G159), .B2(new_n801), .ZN(new_n1093));
  AND4_X1   g0893(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT112), .B(G322), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n801), .A2(new_n1095), .B1(new_n788), .B2(G311), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n514), .B2(new_n796), .C1(new_n1003), .C2(new_n794), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT48), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n858), .B2(new_n804), .C1(new_n538), .C2(new_n799), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT49), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n272), .B1(new_n784), .B2(new_n800), .C1(new_n505), .C2(new_n780), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1094), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1085), .B1(new_n709), .B2(new_n1086), .C1(new_n1104), .C2(new_n841), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT113), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n764), .B2(new_n1040), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1075), .A2(new_n1107), .ZN(G393));
  NOR2_X1   g0908(.A1(new_n1044), .A2(new_n712), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1036), .A2(new_n713), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n764), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n817), .B1(new_n240), .B2(new_n225), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n244), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n821), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n766), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n802), .A2(new_n1003), .B1(new_n794), .B2(new_n856), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n789), .A2(new_n514), .B1(new_n858), .B2(new_n799), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n272), .B1(new_n804), .B2(new_n505), .C1(new_n238), .C2(new_n780), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1095), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1121), .A2(new_n784), .B1(new_n538), .B2(new_n796), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n802), .A2(new_n845), .B1(new_n794), .B2(new_n334), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT51), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n805), .A2(G77), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n263), .C1(new_n601), .C2(new_n780), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n789), .A2(new_n207), .B1(new_n432), .B2(new_n796), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n799), .A2(new_n202), .B1(new_n784), .B2(new_n846), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1118), .A2(new_n1123), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1116), .B1(new_n841), .B2(new_n1131), .C1(new_n1051), .C2(new_n1086), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT107), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(new_n761), .A3(new_n1040), .A4(new_n1037), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1074), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n717), .B1(new_n1137), .B2(new_n1111), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1112), .B(new_n1132), .C1(new_n1136), .C2(new_n1138), .ZN(G390));
  NAND3_X1  g0939(.A1(new_n951), .A2(new_n446), .A3(G330), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT116), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT116), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n951), .A2(new_n446), .A3(new_n1142), .A4(G330), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n984), .A3(new_n639), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n975), .A2(new_n830), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n918), .B1(new_n760), .B2(new_n832), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n920), .A2(new_n703), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n916), .A2(KEYINPUT115), .A3(new_n917), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT115), .B1(new_n916), .B2(new_n917), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n832), .C1(new_n756), .C2(new_n919), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT117), .B1(new_n1157), .B2(new_n1152), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n736), .A2(new_n705), .A3(new_n829), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n956), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n760), .A2(new_n832), .A3(new_n918), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1152), .B1(new_n1159), .B2(new_n956), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n963), .A2(new_n964), .A3(new_n904), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n961), .B(KEYINPUT114), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n961), .B1(new_n1146), .B2(new_n918), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1161), .C1(new_n1168), .C2(new_n970), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n967), .B(new_n966), .C1(new_n976), .C2(new_n961), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1170), .A2(new_n1167), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1148), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1163), .B(new_n1169), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1145), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1162), .A2(new_n1149), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1169), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1172), .B1(new_n1170), .B2(new_n1167), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(new_n717), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n966), .A2(new_n770), .A3(new_n967), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n789), .A2(new_n1011), .B1(new_n780), .B2(new_n207), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n272), .B(new_n1183), .C1(G125), .C2(new_n785), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n805), .A2(G159), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n799), .A2(new_n845), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT54), .B(G143), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1190), .A2(new_n796), .B1(new_n852), .B2(new_n794), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G128), .B2(new_n801), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1184), .A2(new_n1185), .A3(new_n1188), .A4(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n780), .A2(new_n202), .B1(new_n784), .B2(new_n538), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n263), .B(new_n1194), .C1(G87), .C2(new_n807), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G116), .A2(new_n795), .B1(new_n788), .B2(G107), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G97), .A2(new_n797), .B1(new_n801), .B2(G283), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n1126), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n841), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n765), .B1(new_n842), .B2(new_n292), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT118), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1181), .A2(new_n764), .B1(new_n1182), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1180), .A2(new_n1203), .ZN(G378));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n310), .A2(new_n312), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n882), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n632), .A2(new_n306), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n323), .A2(new_n1206), .A3(new_n882), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n947), .B2(new_n703), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n911), .B1(new_n1165), .B2(new_n922), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1215), .B(G330), .C1(new_n1218), .C2(new_n921), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n979), .A2(new_n1217), .A3(new_n969), .A4(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1217), .A2(new_n1219), .B1(new_n969), .B2(new_n979), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1205), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n980), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1217), .A2(new_n969), .A3(new_n979), .A4(new_n1219), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(KEYINPUT122), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1224), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1145), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n717), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1222), .A2(new_n764), .A3(new_n1226), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n765), .B1(new_n842), .B2(G50), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n789), .A2(new_n240), .B1(new_n784), .B2(new_n858), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n272), .A2(new_n478), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1088), .A3(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n795), .A2(KEYINPUT121), .A3(G107), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT121), .B1(new_n795), .B2(G107), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1015), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n780), .A2(new_n201), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n796), .A2(new_n435), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(G116), .C2(new_n801), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1240), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT58), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1239), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT120), .Z(new_n1251));
  AND2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n789), .A2(new_n852), .B1(new_n1253), .B2(new_n794), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n801), .A2(G125), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n1011), .B2(new_n796), .C1(new_n799), .C2(new_n1190), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G150), .C2(new_n805), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT59), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n781), .A2(G159), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1252), .B1(new_n1248), .B2(new_n1247), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1237), .B1(new_n1264), .B2(new_n777), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1215), .B2(new_n771), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1236), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1235), .A2(new_n1268), .ZN(G375));
  NAND3_X1  g1069(.A1(new_n1145), .A2(new_n1149), .A3(new_n1162), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1176), .A2(new_n1049), .A3(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G132), .A2(new_n801), .B1(new_n788), .B2(new_n1189), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1011), .B2(new_n794), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT124), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n799), .A2(new_n334), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n796), .A2(new_n845), .B1(new_n784), .B2(new_n1253), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n263), .B1(new_n804), .B2(new_n207), .C1(new_n201), .C2(new_n780), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(KEYINPUT124), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n272), .B1(new_n780), .B2(new_n383), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT123), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1087), .B1(new_n858), .B2(new_n794), .C1(new_n789), .C2(new_n505), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n802), .A2(new_n538), .B1(new_n799), .B2(new_n240), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n796), .A2(new_n238), .B1(new_n784), .B2(new_n514), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1278), .A2(new_n1279), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n765), .B1(G68), .B2(new_n842), .C1(new_n1286), .C2(new_n841), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1153), .B2(new_n770), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1175), .B2(new_n764), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1271), .A2(new_n1289), .ZN(G381));
  AOI21_X1  g1090(.A(new_n1233), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1267), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1180), .A3(new_n1203), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  INV_X1    g1095(.A(G396), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1075), .A2(new_n1296), .A3(new_n1107), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  OR4_X1    g1099(.A1(G387), .A2(new_n1293), .A3(G381), .A4(new_n1299), .ZN(G407));
  OAI211_X1 g1100(.A(G407), .B(G213), .C1(G343), .C2(new_n1293), .ZN(G409));
  OAI21_X1  g1101(.A(G378), .B1(new_n1291), .B2(new_n1267), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1224), .A2(new_n764), .A3(new_n1225), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1180), .A2(new_n1203), .A3(new_n1266), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1222), .A2(new_n1049), .A3(new_n1227), .A4(new_n1226), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1305), .A2(new_n1306), .B1(G213), .B2(new_n697), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1270), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1149), .A4(new_n1162), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1176), .A3(new_n717), .A4(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(G384), .A3(new_n1289), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1311), .B2(new_n1289), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1302), .A2(new_n1307), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1302), .A2(new_n1307), .A3(KEYINPUT63), .A4(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1062), .B(new_n1064), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1049), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1135), .B2(new_n761), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1324), .B2(new_n764), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1069), .B1(new_n1325), .B2(new_n1024), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1070), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1294), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1067), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1296), .B1(new_n1075), .B2(new_n1107), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1298), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1331), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(KEYINPUT125), .A3(new_n1297), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1329), .A2(G390), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1328), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(G390), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1325), .A2(new_n1024), .A3(G390), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(KEYINPUT126), .B1(new_n1338), .B2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1329), .A2(G390), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1340), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1332), .B(new_n1334), .C1(new_n1343), .C2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1337), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n697), .A2(G213), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1306), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1347), .B1(new_n1348), .B2(new_n1304), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(G375), .B2(G378), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1314), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n697), .A2(G213), .A3(G2897), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n1312), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1352), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1321), .B(new_n1346), .C1(new_n1350), .C2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(KEYINPUT127), .B1(new_n1320), .B2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1356), .B1(new_n1302), .B2(new_n1307), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1337), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1359), .A2(new_n1360), .A3(KEYINPUT61), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1361), .A2(new_n1362), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1358), .A2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1359), .A2(KEYINPUT61), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1360), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1364), .A2(new_n1369), .ZN(G405));
  AND2_X1   g1170(.A1(new_n1293), .A2(new_n1302), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1315), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1373), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1346), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  OR2_X1    g1176(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1377), .A2(new_n1360), .A3(new_n1373), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1376), .A2(new_n1378), .ZN(G402));
endmodule


