//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT64), .A2(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n191), .A2(new_n192), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n189), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT64), .A2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G143), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(G128), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n198), .B1(new_n191), .B2(new_n192), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n189), .A2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n197), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G104), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(G107), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n221), .B1(new_n214), .B2(new_n216), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(KEYINPUT80), .A3(new_n219), .A4(new_n218), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n219), .B1(new_n216), .B2(new_n221), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n231), .A2(KEYINPUT84), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT84), .B1(new_n231), .B2(new_n235), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT10), .B(new_n213), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n227), .A2(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n195), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n194), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n210), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n243), .B2(new_n200), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(KEYINPUT82), .C1(new_n199), .C2(new_n190), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n194), .A2(new_n196), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n223), .B1(new_n222), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(G101), .B1(new_n228), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT64), .B(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n243), .B1(new_n254), .B2(new_n198), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G128), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT65), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n194), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(G101), .C1(new_n228), .C2(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n211), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND4_X1   g078(.A1(new_n257), .A2(new_n259), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n248), .A2(new_n249), .B1(new_n253), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT66), .B(G131), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(new_n269), .A3(new_n271), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n238), .A2(new_n266), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G227), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  INV_X1    g100(.A(new_n248), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n236), .A2(new_n237), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n212), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n286), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n231), .A2(new_n235), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n239), .A2(KEYINPUT84), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n212), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n278), .B1(new_n295), .B2(new_n248), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n285), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n278), .B1(new_n238), .B2(new_n266), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n284), .B1(new_n300), .B2(new_n279), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n187), .B(new_n188), .C1(new_n298), .C2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n284), .A3(new_n279), .ZN(new_n303));
  INV_X1    g117(.A(new_n279), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n290), .B2(new_n297), .ZN(new_n305));
  OAI211_X1 g119(.A(G469), .B(new_n303), .C1(new_n305), .C2(new_n284), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n187), .A2(new_n188), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT77), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT78), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G952), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(G234), .B2(G237), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n188), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT21), .B(G898), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT2), .B(G113), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G116), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n328), .A3(G119), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT69), .B1(new_n325), .B2(G119), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT68), .B(G116), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G119), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n330), .B1(new_n333), .B2(G119), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT5), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G116), .ZN(new_n341));
  OAI21_X1  g155(.A(G113), .B1(new_n341), .B2(KEYINPUT5), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n336), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n236), .B2(new_n237), .ZN(new_n345));
  XNOR2_X1  g159(.A(G110), .B(G122), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n347));
  INV_X1    g161(.A(new_n324), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n337), .B2(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n332), .A2(new_n335), .A3(new_n324), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n219), .B1(new_n229), .B2(new_n218), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n260), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n253), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n227), .B2(new_n230), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n332), .A2(new_n335), .A3(new_n324), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n261), .B1(new_n356), .B2(new_n336), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT85), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n345), .A2(new_n346), .A3(new_n353), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n256), .B1(new_n209), .B2(new_n210), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n360), .A2(new_n262), .B1(new_n194), .B2(new_n258), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G125), .A3(new_n257), .ZN(new_n362));
  INV_X1    g176(.A(G224), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT87), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(new_n365), .C1(new_n212), .C2(G125), .ZN(new_n366));
  INV_X1    g180(.A(new_n364), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT86), .B1(new_n239), .B2(new_n344), .ZN(new_n371));
  INV_X1    g185(.A(new_n344), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n291), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n345), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n346), .B(KEYINPUT8), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n375), .A2(new_n376), .B1(new_n366), .B2(new_n368), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n346), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n358), .A2(new_n353), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n372), .B1(new_n293), .B2(new_n294), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n362), .B1(new_n212), .B2(G125), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(new_n367), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n378), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n378), .B2(new_n388), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n322), .B(new_n323), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n220), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n316), .A3(G214), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(G143), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT88), .B1(new_n397), .B2(new_n275), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n198), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n400));
  INV_X1    g214(.A(new_n275), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n275), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G125), .ZN(new_n406));
  INV_X1    g220(.A(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT16), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n407), .A2(KEYINPUT16), .A3(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G146), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n406), .A2(new_n408), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(KEYINPUT89), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n414), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n404), .B(new_n411), .C1(new_n254), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n418));
  INV_X1    g232(.A(G131), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n397), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n399), .A2(KEYINPUT18), .A3(G131), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n193), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n189), .B2(new_n412), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n394), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n427), .A2(new_n398), .A3(new_n402), .A4(new_n403), .ZN(new_n428));
  INV_X1    g242(.A(new_n411), .ZN(new_n429));
  AOI21_X1  g243(.A(G146), .B1(new_n409), .B2(new_n410), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n398), .A2(new_n402), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(KEYINPUT17), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n428), .B1(new_n433), .B2(KEYINPUT90), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n427), .B1(new_n398), .B2(new_n402), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(new_n431), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n426), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n425), .B1(new_n438), .B2(new_n394), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT20), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n433), .A2(KEYINPUT90), .ZN(new_n443));
  INV_X1    g257(.A(new_n428), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n437), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n394), .A3(new_n424), .ZN(new_n446));
  INV_X1    g260(.A(new_n425), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n440), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n394), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n452), .B(new_n426), .C1(new_n434), .C2(new_n437), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n394), .B1(new_n445), .B2(new_n424), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n188), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G475), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n311), .A2(new_n457), .A3(G953), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n333), .A2(G122), .ZN(new_n459));
  AND2_X1   g273(.A1(KEYINPUT91), .A2(G122), .ZN(new_n460));
  NOR2_X1   g274(.A1(KEYINPUT91), .A2(G122), .ZN(new_n461));
  OAI21_X1  g275(.A(G116), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G107), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n462), .A3(new_n215), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G128), .B(G143), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT13), .B1(new_n195), .B2(G143), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n268), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n467), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n459), .B2(KEYINPUT14), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n333), .A2(KEYINPUT92), .A3(new_n474), .A4(G122), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(KEYINPUT14), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n462), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n477), .A2(G107), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n467), .A2(G134), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n467), .A2(G134), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n458), .B(new_n471), .C1(new_n478), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n458), .ZN(new_n483));
  INV_X1    g297(.A(new_n471), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n477), .B2(G107), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT93), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n188), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n490), .B(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n451), .A2(new_n456), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n315), .A2(new_n392), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n457), .B1(G234), .B2(new_n188), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n340), .A2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n340), .A2(G128), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(KEYINPUT23), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  XNOR2_X1  g317(.A(G119), .B(G128), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(G110), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n429), .B2(new_n430), .ZN(new_n506));
  OAI22_X1  g320(.A1(new_n502), .A2(G110), .B1(new_n503), .B2(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n411), .A3(new_n422), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(G221), .A2(G234), .ZN(new_n510));
  OR3_X1    g324(.A1(new_n510), .A2(KEYINPUT74), .A3(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT74), .B1(new_n510), .B2(G953), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT25), .B1(new_n520), .B2(new_n188), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n516), .B1(new_n506), .B2(new_n508), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT25), .B(new_n188), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n498), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n528), .B(new_n498), .C1(new_n521), .C2(new_n525), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n498), .A2(G902), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  INV_X1    g349(.A(new_n276), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n270), .A2(G134), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n419), .B1(new_n537), .B2(new_n272), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n195), .B1(new_n540), .B2(KEYINPUT67), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n255), .B1(new_n541), .B2(new_n207), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(new_n197), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n257), .A2(new_n277), .A3(new_n259), .A4(new_n264), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n361), .A2(new_n546), .A3(new_n277), .A4(new_n257), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n356), .B2(new_n336), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n349), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n543), .A2(new_n552), .A3(new_n545), .A4(new_n547), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n535), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n539), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n544), .B1(new_n212), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT28), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n395), .A2(new_n316), .A3(G210), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT27), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT26), .B(G101), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(KEYINPUT29), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n188), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n349), .A2(new_n350), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n558), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n535), .B1(new_n570), .B2(new_n555), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n565), .B1(new_n571), .B2(new_n560), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n558), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n543), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n547), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n569), .ZN(new_n576));
  INV_X1    g390(.A(new_n565), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n555), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT29), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G472), .B1(new_n568), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n574), .A2(new_n575), .A3(new_n569), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n555), .A2(new_n565), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT31), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n577), .B1(new_n571), .B2(new_n560), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n576), .A2(new_n585), .A3(new_n555), .A4(new_n565), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT72), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n594), .B(KEYINPUT32), .C1(new_n587), .C2(new_n588), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n596));
  NOR4_X1   g410(.A1(new_n590), .A2(new_n593), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n593), .A2(new_n595), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n599));
  INV_X1    g413(.A(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n561), .B2(new_n566), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(G472), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT73), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n497), .B(new_n534), .C1(new_n597), .C2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  INV_X1    g420(.A(new_n392), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n285), .A2(new_n299), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n286), .B(new_n278), .C1(new_n295), .C2(new_n248), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n279), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n611), .B2(new_n283), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n307), .B1(new_n612), .B2(G469), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n313), .B1(new_n613), .B2(new_n302), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n587), .A2(new_n188), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n534), .A2(new_n616), .A3(new_n591), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n607), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n451), .A2(new_n456), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n488), .A2(new_n620), .A3(new_n489), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n482), .A2(new_n486), .A3(KEYINPUT33), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(G478), .A3(new_n188), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n490), .A2(new_n491), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT94), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AOI211_X1 g445(.A(KEYINPUT20), .B(new_n441), .C1(new_n446), .C2(new_n447), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(KEYINPUT95), .B1(new_n455), .B2(G475), .ZN(new_n633));
  INV_X1    g447(.A(new_n494), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n442), .A2(new_n450), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n509), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n532), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n527), .A2(new_n529), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n527), .A2(KEYINPUT96), .A3(new_n529), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n591), .A3(new_n616), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n607), .A2(new_n650), .A3(new_n614), .A4(new_n495), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT97), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G12));
  NAND2_X1  g468(.A1(new_n591), .A2(new_n592), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n594), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT32), .B1(new_n587), .B2(new_n588), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT72), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n596), .B1(new_n659), .B2(new_n590), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n598), .A2(new_n603), .A3(KEYINPUT73), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n318), .B1(new_n319), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n378), .A2(new_n388), .ZN(new_n668));
  INV_X1    g482(.A(new_n389), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n378), .A2(new_n388), .A3(new_n389), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n672), .A3(KEYINPUT98), .A4(new_n323), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n323), .B1(new_n390), .B2(new_n391), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(new_n666), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n662), .A2(new_n677), .A3(new_n614), .A4(new_n649), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NAND3_X1  g493(.A1(new_n554), .A2(new_n555), .A3(new_n577), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n188), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n577), .B1(new_n576), .B2(new_n555), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n589), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n656), .A2(new_n684), .A3(new_n658), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n598), .A2(KEYINPUT99), .A3(new_n684), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n672), .B(KEYINPUT38), .Z(new_n690));
  INV_X1    g504(.A(new_n649), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n323), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n494), .B1(new_n451), .B2(new_n456), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n690), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n664), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n614), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n689), .A2(new_n698), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n198), .ZN(G45));
  NOR3_X1   g518(.A1(new_n619), .A2(new_n626), .A3(new_n664), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n675), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n662), .A2(new_n614), .A3(new_n707), .A4(new_n649), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n534), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n660), .B2(new_n661), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n188), .B1(new_n298), .B2(new_n301), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n314), .A3(new_n302), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n607), .A2(new_n627), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NOR2_X1   g534(.A1(new_n392), .A2(new_n637), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT101), .B(G116), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G18));
  NAND2_X1  g538(.A1(new_n495), .A2(new_n322), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n714), .A3(new_n675), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n649), .B(new_n726), .C1(new_n597), .C2(new_n604), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR2_X1   g542(.A1(new_n714), .A2(new_n675), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n577), .B1(new_n556), .B2(new_n560), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n583), .A3(new_n586), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n588), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n588), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n534), .A2(new_n734), .A3(new_n616), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n694), .A2(new_n321), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n729), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  AND4_X1   g553(.A1(new_n616), .A2(new_n734), .A3(new_n649), .A4(new_n735), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n705), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n675), .A3(new_n714), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n407), .ZN(G27));
  NAND3_X1  g557(.A1(new_n670), .A2(new_n323), .A3(new_n671), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n315), .A2(new_n710), .A3(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n705), .B(new_n745), .C1(new_n597), .C2(new_n604), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n662), .A2(KEYINPUT103), .A3(new_n705), .A4(new_n745), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n599), .B2(new_n657), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n655), .A2(KEYINPUT105), .A3(new_n589), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n580), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n745), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(KEYINPUT106), .A3(new_n745), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT107), .B1(new_n751), .B2(new_n761), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  OAI211_X1 g580(.A(new_n667), .B(new_n745), .C1(new_n597), .C2(new_n604), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT108), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n662), .A2(new_n769), .A3(new_n667), .A4(new_n745), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n619), .A2(new_n625), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n619), .A2(new_n775), .A3(new_n625), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n616), .A2(new_n591), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n649), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n670), .A2(new_n323), .A3(new_n671), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n777), .B2(new_n779), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(G469), .B1(new_n612), .B2(KEYINPUT45), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n786), .B(new_n608), .C1(new_n611), .C2(new_n283), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n308), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n302), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n313), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n699), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n784), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  OR2_X1    g610(.A1(new_n793), .A2(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n662), .A2(new_n534), .A3(new_n706), .A4(new_n744), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NAND2_X1  g616(.A1(new_n614), .A2(new_n782), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n741), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n768), .B2(new_n770), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n625), .B1(new_n451), .B2(new_n456), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n495), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n607), .A2(new_n614), .A3(new_n807), .A4(new_n617), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n738), .A2(new_n651), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n605), .A3(new_n727), .ZN(new_n810));
  INV_X1    g624(.A(new_n717), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n711), .B(new_n715), .C1(new_n811), .C2(new_n721), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n633), .A2(new_n636), .A3(new_n494), .A4(new_n665), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n315), .A2(new_n813), .A3(new_n744), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n649), .B(new_n814), .C1(new_n597), .C2(new_n604), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n662), .A2(KEYINPUT111), .A3(new_n649), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n805), .A2(new_n810), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n763), .A2(new_n820), .A3(new_n764), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  INV_X1    g636(.A(new_n742), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n678), .A2(new_n823), .A3(new_n708), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n672), .A2(new_n323), .A3(new_n693), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n645), .A2(new_n664), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n309), .A2(new_n314), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT99), .B1(new_n598), .B2(new_n684), .ZN(new_n830));
  AND4_X1   g644(.A1(KEYINPUT99), .A2(new_n656), .A3(new_n658), .A4(new_n684), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n825), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n825), .B1(new_n689), .B2(new_n829), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n822), .B1(new_n824), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n822), .B(new_n837), .C1(new_n824), .C2(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n821), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n750), .B1(new_n746), .B2(new_n747), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n614), .A2(new_n534), .A3(new_n782), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n660), .B2(new_n661), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT103), .B1(new_n845), .B2(new_n705), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n761), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT107), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n804), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n771), .A2(new_n819), .A3(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n605), .A2(new_n812), .A3(new_n727), .A4(new_n809), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n851), .A3(new_n762), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n824), .B2(new_n835), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n315), .B(new_n691), .C1(new_n660), .C2(new_n661), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n742), .B1(new_n856), .B2(new_n677), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n832), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n708), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n863));
  NOR3_X1   g677(.A1(new_n853), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n842), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n853), .B2(new_n862), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n820), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n841), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n714), .A2(new_n323), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT116), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n318), .A2(new_n736), .A3(new_n774), .A4(new_n776), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n690), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n873), .A2(KEYINPUT50), .A3(new_n874), .A4(new_n690), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n714), .A2(new_n744), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n318), .A2(new_n880), .A3(new_n774), .A4(new_n776), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n740), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n881), .B2(new_n740), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n689), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n880), .A2(new_n534), .A3(new_n318), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n619), .A3(new_n626), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n879), .A2(new_n885), .A3(KEYINPUT51), .A4(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n713), .A2(new_n302), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n797), .B(new_n798), .C1(new_n314), .C2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n874), .A2(new_n782), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n892), .B2(KEYINPUT118), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n879), .A2(new_n885), .A3(new_n888), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n782), .A3(new_n874), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT51), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n881), .A2(new_n534), .A3(new_n756), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n886), .A2(new_n627), .A3(new_n887), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n317), .B(KEYINPUT119), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n874), .B2(new_n729), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n896), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n865), .A2(new_n871), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(G952), .A2(G953), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n891), .A2(KEYINPUT49), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT109), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n534), .A2(new_n314), .A3(new_n323), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n773), .B(new_n912), .C1(new_n891), .C2(KEYINPUT49), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n911), .A2(new_n886), .A3(new_n690), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT110), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n316), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n866), .A2(new_n870), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n188), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n383), .A2(new_n385), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n387), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n922), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT56), .B(new_n928), .C1(new_n924), .C2(G210), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G51));
  NAND2_X1  g746(.A1(new_n866), .A2(new_n870), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n867), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n307), .B(KEYINPUT57), .Z(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n301), .B2(new_n298), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n785), .A2(new_n787), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n921), .B1(new_n936), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n921), .B1(new_n940), .B2(new_n439), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .A4(new_n448), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(G60));
  AND2_X1   g757(.A1(new_n621), .A2(new_n622), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n922), .B1(new_n934), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n865), .B2(new_n871), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G63));
  XNOR2_X1  g766(.A(new_n520), .B(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n923), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n866), .B2(new_n870), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n921), .B1(new_n957), .B2(new_n643), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT122), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT61), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n956), .B(new_n958), .C1(KEYINPUT122), .C2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(G66));
  XOR2_X1   g778(.A(new_n852), .B(KEYINPUT123), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n316), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n320), .B2(new_n363), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n926), .B1(G898), .B2(new_n316), .ZN(new_n969));
  XOR2_X1   g783(.A(KEYINPUT124), .B(KEYINPUT125), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n968), .B(new_n971), .ZN(G69));
  NAND2_X1  g786(.A1(new_n574), .A2(new_n575), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n416), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n703), .A2(KEYINPUT62), .A3(new_n824), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n700), .A2(new_n495), .A3(new_n744), .A4(new_n806), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n784), .A2(new_n794), .B1(new_n711), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT62), .B1(new_n703), .B2(new_n824), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n975), .A2(new_n977), .A3(new_n801), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(new_n316), .ZN(new_n980));
  INV_X1    g794(.A(new_n824), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n756), .A2(new_n534), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n826), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n794), .B1(new_n784), .B2(new_n983), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n771), .A2(new_n801), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n316), .A3(new_n765), .ZN(new_n986));
  INV_X1    g800(.A(new_n974), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(G900), .B2(G953), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n980), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(G953), .B1(new_n281), .B2(new_n663), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G72));
  INV_X1    g805(.A(new_n578), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n992), .A2(new_n682), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n842), .B2(new_n864), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT127), .Z(new_n998));
  OAI21_X1  g812(.A(new_n994), .B1(new_n979), .B2(new_n965), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n921), .B1(new_n999), .B2(new_n682), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n985), .A2(new_n765), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n994), .B1(new_n1001), .B2(new_n965), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n992), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n998), .A2(new_n1006), .ZN(G57));
endmodule


