//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n463), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(new_n463), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n476), .B2(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n473), .A2(new_n474), .A3(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G136), .B2(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n474), .A3(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n473), .A2(new_n463), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n500), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n494), .B1(new_n503), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT6), .B(G651), .Z(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n521), .A3(KEYINPUT70), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT71), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n520), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n509), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n534), .A3(KEYINPUT72), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n524), .B2(new_n525), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(new_n533), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n535), .A2(new_n540), .ZN(G168));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n526), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n509), .A2(new_n520), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n544), .A2(new_n511), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n551), .A2(new_n511), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n526), .B2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  AND2_X1   g134(.A1(new_n518), .A2(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(KEYINPUT74), .A3(new_n511), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT74), .B1(new_n563), .B2(new_n511), .ZN(new_n565));
  INV_X1    g140(.A(new_n545), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n543), .A2(new_n570), .A3(new_n548), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND2_X1  g150(.A1(new_n566), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n522), .C2(new_n578), .ZN(G288));
  AND2_X1   g154(.A1(G48), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n520), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n511), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n545), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n583), .A2(new_n585), .ZN(G305));
  AND2_X1   g161(.A1(new_n526), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n511), .B1(new_n545), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n526), .A2(G54), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n545), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n532), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n594), .A2(new_n597), .B1(G651), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n572), .B2(G868), .ZN(G284));
  AOI21_X1  g179(.A(new_n603), .B1(new_n572), .B2(G868), .ZN(G321));
  NOR2_X1   g180(.A1(G299), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g182(.A(new_n606), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(new_n602), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  INV_X1    g186(.A(new_n554), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n602), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n477), .A2(new_n499), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n504), .A2(new_n474), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n489), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n474), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n621), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT77), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  NOR2_X1   g221(.A1(G2072), .A2(G2078), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n442), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT17), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT78), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT80), .Z(new_n654));
  OR2_X1    g229(.A1(new_n648), .A2(KEYINPUT79), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n648), .A2(KEYINPUT79), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n652), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n649), .C2(new_n651), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n651), .A2(new_n648), .A3(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n673), .S(new_n666), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT81), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(new_n687), .ZN(G229));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT86), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NOR2_X1   g270(.A1(G166), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G22), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(G288), .A2(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G23), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT87), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n699), .B(new_n700), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n706), .B2(new_n704), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n693), .A2(new_n694), .A3(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n591), .A2(new_n695), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n695), .B2(G24), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(new_n686), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT85), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n489), .A2(G131), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n622), .A2(G119), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n713), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G1986), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n710), .A2(new_n711), .A3(new_n714), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT36), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n488), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT89), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(new_n474), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G33), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  OAI21_X1  g314(.A(KEYINPUT90), .B1(G29), .B2(G32), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n622), .A2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n489), .A2(G141), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n477), .A2(G105), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(KEYINPUT90), .B(new_n740), .S(new_n750), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  INV_X1    g329(.A(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT24), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n479), .B2(new_n749), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n739), .B(new_n753), .C1(new_n754), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n609), .A2(new_n695), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G4), .B2(new_n695), .ZN(new_n762));
  INV_X1    g337(.A(G1348), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n752), .B2(new_n751), .ZN(new_n765));
  NAND2_X1  g340(.A1(G164), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G27), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n749), .B1(new_n772), .B2(G28), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(G28), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(KEYINPUT92), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n771), .B1(new_n774), .B2(new_n776), .C1(new_n627), .C2(new_n749), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n765), .A2(new_n769), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n695), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n554), .B2(new_n695), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1341), .ZN(new_n781));
  NOR2_X1   g356(.A1(G29), .A2(G35), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G162), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2090), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n695), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n695), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n762), .A2(new_n763), .B1(new_n790), .B2(G1961), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n795));
  INV_X1    g370(.A(G140), .ZN(new_n796));
  INV_X1    g371(.A(G128), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n795), .B1(new_n796), .B2(new_n488), .C1(new_n485), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n749), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n758), .A2(new_n754), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n793), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n778), .A2(new_n788), .A3(new_n792), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n695), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G299), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT97), .B(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n786), .B2(new_n787), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G21), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G168), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1966), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n807), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n760), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n728), .A2(new_n820), .ZN(G311));
  INV_X1    g396(.A(G311), .ZN(G150));
  NAND2_X1  g397(.A1(new_n566), .A2(G93), .ZN(new_n823));
  INV_X1    g398(.A(new_n525), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT70), .B1(new_n518), .B2(new_n521), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  OAI211_X1 g402(.A(KEYINPUT99), .B(new_n823), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n827), .B1(new_n524), .B2(new_n525), .ZN(new_n830));
  INV_X1    g405(.A(new_n823), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n511), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n609), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n612), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n833), .A2(new_n554), .A3(new_n835), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n845), .B2(new_n846), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n839), .B1(new_n848), .B2(new_n850), .ZN(G145));
  XOR2_X1   g426(.A(new_n748), .B(new_n798), .Z(new_n852));
  AOI21_X1  g427(.A(new_n495), .B1(new_n484), .B2(new_n505), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT68), .B1(new_n466), .B2(new_n496), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n499), .A2(new_n498), .A3(new_n501), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n491), .B(new_n493), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(G164), .A2(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n861), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n737), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n734), .A2(KEYINPUT103), .A3(new_n736), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n720), .B(new_n619), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n622), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n474), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G142), .B2(new_n489), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n869), .B(new_n874), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n868), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n627), .B(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g456(.A(new_n844), .B(new_n615), .ZN(new_n882));
  XNOR2_X1  g457(.A(G299), .B(new_n602), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n591), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(G303), .B(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n892), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n888), .B(new_n894), .C1(new_n893), .C2(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n613), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n836), .A2(new_n613), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n900), .A2(KEYINPUT105), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n900), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G331));
  INV_X1    g482(.A(new_n843), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n554), .B1(new_n833), .B2(new_n835), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT106), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n842), .B2(new_n843), .ZN(new_n912));
  NAND2_X1  g487(.A1(G286), .A2(new_n549), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n572), .A2(G168), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n908), .B2(new_n909), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n842), .A2(new_n911), .A3(new_n843), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n886), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n915), .B1(new_n910), .B2(new_n912), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n917), .A3(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n884), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(new_n896), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n925), .B2(new_n896), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n892), .B(KEYINPUT104), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n921), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n931), .B2(G37), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT43), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n883), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n886), .B2(KEYINPUT108), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n923), .B2(new_n922), .ZN(new_n937));
  INV_X1    g512(.A(new_n924), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n896), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  AND4_X1   g515(.A1(KEYINPUT43), .A2(new_n934), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n929), .B2(new_n932), .ZN(new_n945));
  AND4_X1   g520(.A1(new_n944), .A2(new_n934), .A3(new_n939), .A4(new_n940), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(G397));
  NOR2_X1   g523(.A1(new_n861), .A2(G1384), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n469), .A2(G40), .A3(new_n478), .A4(new_n475), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n949), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT46), .ZN(new_n954));
  INV_X1    g529(.A(G2067), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n798), .B(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n951), .B1(new_n748), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  INV_X1    g535(.A(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n720), .B(new_n723), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT109), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n748), .B(new_n952), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n956), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n951), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n951), .A2(new_n686), .A3(new_n591), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n967), .A2(KEYINPUT127), .B1(KEYINPUT48), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n970), .B(new_n972), .C1(KEYINPUT127), .C2(new_n967), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n966), .A2(new_n723), .A3(new_n720), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n798), .A2(G2067), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n951), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n962), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n960), .A2(new_n961), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n859), .A2(new_n860), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n950), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(new_n768), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n857), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(G164), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1961), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n950), .B1(new_n857), .B2(new_n991), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n950), .B1(new_n857), .B2(new_n981), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(new_n984), .A3(KEYINPUT53), .A4(new_n768), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n987), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n572), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n857), .B2(new_n989), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n950), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n1007), .B2(new_n982), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n996), .A2(new_n997), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT55), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n698), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n990), .A2(new_n993), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n787), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1013), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n1023));
  INV_X1    g598(.A(new_n583), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT112), .B(G86), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n566), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n678), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n583), .A2(G1981), .A3(new_n585), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1023), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  NOR3_X1   g605(.A1(G164), .A2(G1384), .A3(new_n950), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1015), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1023), .B(new_n1033), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n983), .A2(new_n857), .A3(new_n989), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G288), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1031), .A2(new_n1015), .A3(new_n1039), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(KEYINPUT111), .A3(new_n1043), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1041), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1005), .A2(new_n1014), .A3(new_n1022), .A4(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n535), .A2(new_n540), .A3(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n996), .A2(new_n997), .A3(new_n754), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1966), .B1(new_n1001), .B2(new_n984), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  INV_X1    g633(.A(new_n981), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n983), .B1(G164), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1006), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n996), .A2(new_n997), .A3(new_n754), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1015), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT122), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT51), .B(G8), .C1(new_n1065), .C2(G286), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1057), .A2(new_n1064), .B1(new_n1066), .B2(KEYINPUT121), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1050), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1068), .B(KEYINPUT51), .C1(new_n1063), .C2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n1070), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1049), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1052), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1064), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1066), .A2(KEYINPUT121), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1070), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1081), .B2(KEYINPUT62), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT123), .B(new_n1072), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1073), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1073), .B(KEYINPUT124), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1022), .A2(new_n1014), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1055), .A2(G286), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1048), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(KEYINPUT116), .A3(new_n1091), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1055), .A2(new_n1091), .A3(G286), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1048), .A2(KEYINPUT114), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1048), .A2(KEYINPUT114), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1088), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1022), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G288), .A2(G1976), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT115), .Z(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1034), .B2(new_n1030), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1032), .B1(new_n1105), .B2(new_n1028), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n562), .B2(new_n567), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1018), .B2(G1956), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1009), .A2(KEYINPUT117), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1007), .A2(new_n982), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n994), .A2(new_n763), .A3(new_n999), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(G2067), .B2(new_n1036), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n609), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(KEYINPUT119), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT117), .B1(new_n1009), .B2(new_n1114), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1112), .B(G1956), .C1(new_n996), .C2(new_n997), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G299), .B(KEYINPUT57), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT119), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1119), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1119), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1127), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1016), .B2(G1996), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1007), .A2(KEYINPUT120), .A3(new_n952), .A4(new_n982), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1036), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n554), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1121), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1120), .B(KEYINPUT60), .C1(G2067), .C2(new_n1036), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n609), .A3(new_n1147), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1121), .A2(new_n1145), .A3(new_n609), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1130), .B1(new_n1135), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n950), .A2(new_n986), .A3(G2078), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n982), .B(new_n1153), .C1(new_n949), .C2(KEYINPUT45), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1154), .A2(new_n1000), .A3(new_n987), .ZN(new_n1155));
  OAI221_X1 g730(.A(KEYINPUT54), .B1(new_n572), .B2(new_n1003), .C1(new_n1155), .C2(new_n549), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1154), .A2(new_n987), .A3(G301), .A4(new_n1000), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1004), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1048), .A2(new_n1022), .A3(new_n1014), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1081), .A2(new_n1156), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1107), .B1(new_n1152), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1086), .A2(new_n1087), .A3(new_n1100), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(new_n967), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n591), .B(new_n686), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n951), .B2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT110), .Z(new_n1169));
  AND3_X1   g744(.A1(new_n1164), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1165), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n979), .B1(new_n1170), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g747(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1174));
  OAI211_X1 g748(.A(new_n1174), .B(new_n880), .C1(new_n945), .C2(new_n946), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


