//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G57gat), .B(G64gat), .Z(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n202), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT21), .ZN(new_n214));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n214), .B(new_n215), .Z(new_n216));
  XOR2_X1   g015(.A(G127gat), .B(G155gat), .Z(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT20), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n216), .B(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G183gat), .B(G211gat), .Z(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n221), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n227), .B1(new_n226), .B2(new_n229), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(KEYINPUT21), .B2(new_n213), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n236), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n238), .A3(new_n223), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT41), .ZN(new_n243));
  XNOR2_X1  g042(.A(G134gat), .B(G162gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n243), .B(new_n244), .Z(new_n245));
  AND2_X1   g044(.A1(new_n245), .A2(KEYINPUT96), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G85gat), .A2(G92gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT94), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT94), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(G85gat), .A3(G92gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT7), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT7), .ZN(new_n255));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT8), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT95), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  INV_X1    g058(.A(G92gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n257), .B2(new_n261), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n254), .B(new_n255), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G99gat), .B(G106gat), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n255), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT7), .B1(new_n249), .B2(new_n251), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n257), .A2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT95), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n265), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278));
  NOR4_X1   g077(.A1(new_n278), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n280));
  INV_X1    g079(.A(G36gat), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT85), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n277), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT86), .B(new_n277), .C1(new_n279), .C2(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT15), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT83), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(KEYINPUT83), .B1(G43gat), .B2(G50gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT84), .B(G50gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(G43gat), .ZN(new_n291));
  OR2_X1    g090(.A1(G43gat), .A2(G50gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G43gat), .A2(G50gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G29gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n285), .A2(new_n286), .A3(new_n291), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299));
  NOR3_X1   g098(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n300), .A2(KEYINPUT82), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n277), .B1(new_n300), .B2(KEYINPUT82), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n303), .B2(new_n296), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n299), .B1(new_n298), .B2(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n276), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G190gat), .B(G218gat), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n276), .ZN(new_n310));
  INV_X1    g109(.A(new_n277), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(new_n295), .A3(new_n281), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n278), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n280), .A2(KEYINPUT85), .A3(new_n281), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n291), .B(new_n297), .C1(new_n316), .C2(KEYINPUT86), .ZN(new_n317));
  INV_X1    g116(.A(new_n286), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n304), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n310), .A2(new_n319), .B1(KEYINPUT41), .B2(new_n242), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n307), .A2(new_n309), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n309), .B1(new_n307), .B2(new_n320), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n247), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n245), .A2(KEYINPUT96), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n246), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT97), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n264), .B2(new_n265), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n264), .A2(new_n265), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n274), .B1(new_n269), .B2(new_n273), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(new_n213), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n266), .B(new_n275), .C1(new_n333), .C2(new_n212), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT10), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n276), .A2(new_n340), .A3(new_n212), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(G230gat), .A3(G233gat), .A4(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n241), .A2(new_n331), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G169gat), .ZN(new_n356));
  INV_X1    g155(.A(G176gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n358), .A2(KEYINPUT26), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT27), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G183gat), .ZN(new_n367));
  INV_X1    g166(.A(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT66), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT27), .B(G183gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT28), .A3(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT66), .B1(new_n369), .B2(new_n370), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n363), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n361), .A2(new_n381), .B1(G169gat), .B2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n368), .ZN(new_n383));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT24), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n380), .A2(new_n382), .A3(new_n385), .A4(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n392));
  XOR2_X1   g191(.A(G127gat), .B(G134gat), .Z(new_n393));
  XNOR2_X1  g192(.A(G113gat), .B(G120gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n393), .B1(new_n394), .B2(KEYINPUT1), .ZN(new_n395));
  XOR2_X1   g194(.A(G113gat), .B(G120gat), .Z(new_n396));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n376), .A2(new_n401), .A3(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n404), .B(KEYINPUT64), .Z(new_n405));
  AND2_X1   g204(.A1(new_n395), .A2(new_n399), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT67), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G15gat), .B(G43gat), .Z(new_n411));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n405), .B1(new_n403), .B2(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT34), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI211_X1 g216(.A(KEYINPUT34), .B(new_n405), .C1(new_n403), .C2(new_n407), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n415), .A2(new_n416), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n410), .B(new_n413), .C1(new_n423), .C2(new_n418), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n420), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT2), .ZN(new_n430));
  INV_X1    g229(.A(new_n429), .ZN(new_n431));
  NOR2_X1   g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G148gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(G141gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT71), .B(G148gat), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(G141gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G148gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n442), .A3(G141gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n435), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n432), .ZN(new_n447));
  XNOR2_X1  g246(.A(G141gat), .B(G148gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450));
  INV_X1    g249(.A(G141gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(G148gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n435), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n453), .A3(new_n430), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n439), .A2(new_n446), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT22), .ZN(new_n457));
  INV_X1    g256(.A(G211gat), .ZN(new_n458));
  INV_X1    g257(.A(G218gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT77), .ZN(new_n462));
  XOR2_X1   g261(.A(G211gat), .B(G218gat), .Z(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n461), .B(new_n463), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT3), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n455), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n443), .A2(new_n438), .A3(new_n444), .ZN(new_n470));
  INV_X1    g269(.A(new_n433), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n446), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n430), .B1(new_n448), .B2(KEYINPUT70), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n435), .A2(new_n452), .A3(new_n450), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n447), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n466), .B1(new_n476), .B2(new_n465), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n428), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n466), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n468), .B1(new_n479), .B2(KEYINPUT29), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n471), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n428), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(KEYINPUT78), .B2(new_n477), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n477), .A2(KEYINPUT78), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(G22gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n478), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT79), .B1(new_n487), .B2(G22gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(G78gat), .B(G106gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G50gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n493), .B(new_n494), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n491), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n488), .A2(KEYINPUT79), .A3(new_n490), .A4(new_n495), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n427), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n376), .A2(new_n390), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n376), .B2(new_n390), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n479), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n376), .A2(new_n390), .A3(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(new_n375), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n373), .A3(new_n371), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n509), .A2(new_n363), .B1(new_n388), .B2(new_n389), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n507), .B(new_n466), .C1(new_n510), .C2(new_n504), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT68), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n503), .A2(new_n505), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n466), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G8gat), .B(G36gat), .Z(new_n517));
  XOR2_X1   g316(.A(G64gat), .B(G92gat), .Z(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(KEYINPUT69), .Z(new_n521));
  NAND3_X1  g320(.A1(new_n512), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n501), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n512), .B2(new_n515), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT30), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT80), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n522), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT30), .B1(new_n528), .B2(new_n525), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT80), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n520), .A2(new_n501), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n500), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT35), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n483), .A2(KEYINPUT3), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n400), .A3(new_n476), .ZN(new_n538));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT5), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n472), .A2(new_n406), .A3(new_n475), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n472), .A2(new_n406), .A3(KEYINPUT4), .A4(new_n475), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n545), .A2(new_n542), .A3(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n540), .B(new_n541), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n538), .A2(new_n545), .A3(new_n546), .A4(new_n539), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n483), .A2(new_n400), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n543), .ZN(new_n553));
  INV_X1    g352(.A(new_n539), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n541), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n550), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G1gat), .B(G29gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT0), .ZN(new_n560));
  XNOR2_X1  g359(.A(G57gat), .B(G85gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(KEYINPUT6), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n538), .A2(new_n541), .A3(new_n539), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT4), .B1(new_n455), .B2(new_n406), .ZN(new_n566));
  INV_X1    g365(.A(new_n546), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT74), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n542), .A3(new_n546), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n557), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n562), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n562), .B(new_n549), .C1(new_n556), .C2(new_n557), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n564), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n535), .A2(new_n536), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n581), .A3(new_n576), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n573), .B2(new_n562), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n558), .A2(KEYINPUT76), .A3(new_n563), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n580), .A2(new_n582), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n564), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n523), .A2(new_n526), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT35), .B1(new_n589), .B2(new_n500), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n588), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n586), .B2(new_n564), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n499), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n425), .B2(new_n426), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n420), .A2(new_n424), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n421), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n420), .A2(new_n424), .A3(new_n422), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT36), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n553), .A2(new_n554), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n538), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n568), .B2(new_n569), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n606), .B2(new_n539), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n538), .B1(new_n548), .B2(new_n547), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n603), .A3(new_n554), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n609), .A3(new_n562), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n610), .A2(new_n611), .B1(new_n558), .B2(new_n563), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT40), .A4(new_n562), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n527), .A2(new_n612), .A3(new_n532), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n499), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n516), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n521), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n506), .A2(new_n511), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(KEYINPUT37), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n525), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n564), .B(new_n622), .C1(new_n574), .C2(new_n577), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n524), .B1(new_n516), .B2(new_n616), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n624), .A2(new_n625), .B1(new_n616), .B2(new_n516), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n601), .B1(new_n615), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n591), .B1(new_n594), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n319), .A2(KEYINPUT17), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n233), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n319), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(new_n232), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n632), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n232), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n233), .A2(new_n319), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n636), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n232), .B1(new_n305), .B2(new_n306), .ZN(new_n650));
  INV_X1    g449(.A(new_n639), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n233), .B2(new_n319), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(KEYINPUT88), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n642), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT90), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n642), .A2(new_n649), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT87), .ZN(new_n658));
  INV_X1    g457(.A(new_n644), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n635), .A2(new_n659), .A3(new_n637), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n650), .A2(new_n644), .A3(new_n636), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT87), .A3(new_n638), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n655), .A2(new_n657), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G113gat), .B(G141gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G197gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(KEYINPUT12), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT91), .B1(new_n673), .B2(new_n654), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n662), .B2(new_n638), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n635), .A2(new_n641), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(KEYINPUT88), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT91), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n642), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n631), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT92), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n631), .B2(new_n682), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n355), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(KEYINPUT98), .B(new_n355), .C1(new_n684), .C2(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n587), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n695));
  INV_X1    g494(.A(new_n691), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n695), .B(G8gat), .C1(new_n696), .C2(new_n533), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n533), .B1(new_n689), .B2(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT99), .B1(new_n698), .B2(new_n227), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n697), .B(new_n699), .C1(new_n702), .C2(new_n703), .ZN(G1325gat));
  INV_X1    g503(.A(new_n427), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n696), .A2(G15gat), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n601), .B(KEYINPUT100), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n696), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n497), .A2(new_n498), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  OR2_X1    g512(.A1(new_n684), .A2(new_n686), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n240), .A2(new_n330), .A3(new_n353), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT101), .Z(new_n716));
  NAND4_X1  g515(.A1(new_n714), .A2(new_n295), .A3(new_n692), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n589), .A2(new_n720), .A3(new_n710), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT103), .B1(new_n593), .B2(new_n499), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n630), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI211_X1 g524(.A(KEYINPUT104), .B(new_n630), .C1(new_n721), .C2(new_n722), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n591), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT105), .B(new_n591), .C1(new_n725), .C2(new_n726), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n331), .A2(KEYINPUT44), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n631), .A2(new_n330), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n240), .B(KEYINPUT102), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n664), .A2(new_n670), .B1(new_n674), .B2(new_n680), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n737), .A2(new_n738), .A3(new_n352), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n740), .B2(new_n587), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G29gat), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n587), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n718), .B1(new_n742), .B2(new_n743), .ZN(G1328gat));
  NAND4_X1  g543(.A1(new_n714), .A2(new_n281), .A3(new_n534), .A4(new_n716), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT46), .Z(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n740), .B2(new_n533), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1329gat));
  OAI21_X1  g547(.A(G43gat), .B1(new_n740), .B2(new_n601), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n714), .A2(new_n716), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n705), .A2(G43gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n739), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n732), .B2(new_n734), .ZN(new_n755));
  INV_X1    g554(.A(new_n707), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(G43gat), .B1(new_n750), .B2(new_n751), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n758), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n499), .A2(new_n290), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n499), .B(new_n754), .C1(new_n732), .C2(new_n734), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n290), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n740), .A2(KEYINPUT107), .A3(new_n499), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n750), .A2(new_n761), .ZN(new_n768));
  INV_X1    g567(.A(new_n290), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n755), .B2(new_n710), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n760), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(G1331gat));
  NOR4_X1   g571(.A1(new_n240), .A2(new_n682), .A3(new_n330), .A4(new_n353), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n729), .A2(new_n730), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n587), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G57gat), .Z(G1332gat));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n729), .A2(KEYINPUT108), .A3(new_n730), .A4(new_n773), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n533), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT109), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n778), .A2(new_n783), .A3(new_n779), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n786));
  INV_X1    g585(.A(G64gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n784), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1333gat));
  NAND4_X1  g590(.A1(new_n778), .A2(G71gat), .A3(new_n756), .A4(new_n779), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n205), .B1(new_n774), .B2(new_n705), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n710), .A3(new_n779), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n241), .A2(new_n682), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n352), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n732), .B2(new_n734), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n587), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n330), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n727), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n692), .A2(new_n259), .A3(new_n352), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  INV_X1    g609(.A(new_n807), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n533), .A2(G92gat), .A3(new_n353), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT110), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT111), .Z(new_n816));
  AND3_X1   g615(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n260), .B1(new_n800), .B2(new_n534), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n799), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n735), .A2(new_n534), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G92gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n815), .B1(new_n806), .B2(new_n807), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT113), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n818), .A2(new_n828), .A3(new_n825), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n819), .B1(new_n827), .B2(new_n829), .ZN(G1337gat));
  OAI21_X1  g629(.A(G99gat), .B1(new_n801), .B2(new_n707), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n705), .A2(G99gat), .A3(new_n353), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n808), .B2(new_n832), .ZN(G1338gat));
  NOR3_X1   g632(.A1(new_n499), .A2(G106gat), .A3(new_n353), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n812), .A2(new_n813), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(G106gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n800), .B2(new_n710), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839));
  INV_X1    g638(.A(new_n834), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n808), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n837), .B2(new_n841), .ZN(G1339gat));
  NOR2_X1   g641(.A1(new_n354), .A2(new_n682), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n637), .B1(new_n635), .B2(new_n659), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n668), .ZN(new_n847));
  AOI221_X4 g646(.A(new_n847), .B1(new_n329), .B2(new_n324), .C1(new_n674), .C2(new_n680), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n332), .C1(new_n339), .C2(new_n341), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n348), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n853), .A3(new_n348), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n339), .A2(new_n332), .A3(new_n341), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(KEYINPUT54), .A3(new_n342), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n850), .A2(new_n853), .A3(new_n348), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n853), .B1(new_n850), .B2(new_n348), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n857), .B(KEYINPUT55), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n350), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT115), .B1(new_n863), .B2(new_n350), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n848), .B(new_n860), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n342), .A2(KEYINPUT54), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n339), .A2(new_n332), .A3(new_n341), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT55), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n854), .B2(new_n852), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(new_n349), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n350), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n860), .A4(new_n848), .ZN(new_n877));
  INV_X1    g676(.A(new_n847), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n681), .A2(new_n352), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT55), .B1(new_n855), .B2(new_n857), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n873), .B2(new_n874), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n881), .B2(new_n682), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n867), .B(new_n877), .C1(new_n882), .C2(new_n330), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n843), .B1(new_n883), .B2(new_n736), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n587), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n535), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n738), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n353), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT117), .B(G120gat), .Z(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(G1341gat));
  OAI21_X1  g690(.A(G127gat), .B1(new_n886), .B2(new_n736), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n240), .A2(G127gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n886), .B2(new_n893), .ZN(G1342gat));
  AOI211_X1 g693(.A(new_n331), .B(new_n886), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1343gat));
  NAND3_X1  g696(.A1(new_n681), .A2(new_n352), .A3(new_n878), .ZN(new_n898));
  INV_X1    g697(.A(new_n871), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n349), .B1(new_n899), .B2(new_n855), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n860), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(new_n738), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n331), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n867), .A3(new_n877), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n843), .B1(new_n904), .B2(new_n240), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n499), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n867), .A2(new_n877), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n682), .B(new_n860), .C1(new_n864), .C2(new_n865), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n330), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n736), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n355), .A2(new_n738), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n710), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n692), .A2(new_n533), .A3(new_n601), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n906), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G141gat), .B1(new_n916), .B2(new_n738), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT58), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n756), .A2(new_n499), .A3(new_n534), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n885), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n682), .A2(new_n451), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n919), .B(new_n923), .Z(G1344gat));
  INV_X1    g723(.A(new_n921), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n436), .A3(new_n352), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT119), .Z(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n499), .A2(KEYINPUT57), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n682), .A2(new_n860), .A3(new_n900), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n330), .B1(new_n932), .B2(new_n898), .ZN(new_n933));
  INV_X1    g732(.A(new_n866), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n880), .A2(new_n872), .A3(new_n349), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n879), .B1(new_n936), .B2(new_n682), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT120), .B(new_n866), .C1(new_n937), .C2(new_n330), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n240), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n930), .B1(new_n939), .B2(new_n911), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n912), .A2(new_n710), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(KEYINPUT57), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n352), .A3(new_n915), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n928), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  INV_X1    g743(.A(new_n916), .ZN(new_n945));
  AOI211_X1 g744(.A(KEYINPUT59), .B(new_n436), .C1(new_n945), .C2(new_n352), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n927), .B1(new_n944), .B2(new_n946), .ZN(G1345gat));
  OR3_X1    g746(.A1(new_n921), .A2(G155gat), .A3(new_n240), .ZN(new_n948));
  OAI21_X1  g747(.A(G155gat), .B1(new_n916), .B2(new_n736), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1346gat));
  AOI21_X1  g749(.A(G162gat), .B1(new_n925), .B2(new_n330), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n330), .A2(G162gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n945), .B2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n884), .A2(new_n692), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n954), .A2(new_n499), .A3(new_n534), .A4(new_n427), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n682), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n692), .A2(new_n533), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT121), .B1(new_n958), .B2(new_n427), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(KEYINPUT121), .A3(new_n427), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n499), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n884), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n738), .A2(new_n356), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n956), .A2(new_n357), .A3(new_n352), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n962), .A2(new_n352), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n357), .ZN(G1349gat));
  AOI21_X1  g766(.A(new_n364), .B1(new_n962), .B2(new_n737), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n241), .A2(new_n372), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n956), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g770(.A(new_n368), .B1(new_n962), .B2(new_n330), .ZN(new_n972));
  XNOR2_X1  g771(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n368), .A3(new_n330), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1351gat));
  NAND3_X1  g775(.A1(new_n707), .A2(new_n710), .A3(new_n534), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT123), .Z(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n954), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(KEYINPUT124), .B(G197gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n682), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n707), .A2(new_n958), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n942), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n985), .A2(new_n738), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n986), .B2(new_n981), .ZN(G1352gat));
  NOR3_X1   g786(.A1(new_n979), .A2(G204gat), .A3(new_n353), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  OAI21_X1  g788(.A(G204gat), .B1(new_n985), .B2(new_n353), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n980), .A2(new_n458), .A3(new_n241), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n913), .B1(new_n912), .B2(new_n710), .ZN(new_n993));
  NOR4_X1   g792(.A1(new_n993), .A2(new_n940), .A3(new_n240), .A4(new_n983), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n458), .B1(new_n994), .B2(KEYINPUT125), .ZN(new_n995));
  OAI21_X1  g794(.A(KEYINPUT57), .B1(new_n884), .B2(new_n499), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n938), .A2(new_n240), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT120), .B1(new_n903), .B2(new_n866), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n911), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(new_n929), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n996), .A2(new_n241), .A3(new_n1000), .A4(new_n984), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n241), .A4(new_n984), .ZN(new_n1005));
  AND4_X1   g804(.A1(KEYINPUT63), .A2(new_n1005), .A3(new_n1003), .A4(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n992), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1009));
  OAI211_X1 g808(.A(new_n1009), .B(new_n992), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(G1354gat));
  AOI21_X1  g810(.A(G218gat), .B1(new_n980), .B2(new_n330), .ZN(new_n1012));
  INV_X1    g811(.A(new_n985), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n330), .A2(G218gat), .ZN(new_n1014));
  XOR2_X1   g813(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  AOI21_X1  g814(.A(new_n1012), .B1(new_n1013), .B2(new_n1015), .ZN(G1355gat));
endmodule


