//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  OR2_X1    g004(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n204), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(G141gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n214), .B(KEYINPUT76), .C1(G141gat), .C2(new_n209), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT77), .A3(new_n216), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n215), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n216), .B(new_n224), .C1(new_n228), .C2(KEYINPUT2), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n203), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232));
  INV_X1    g031(.A(G127gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(G113gat), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G113gat), .B2(G120gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n234), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n241), .B(new_n234), .C1(new_n237), .C2(new_n239), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n203), .A3(new_n229), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n245), .A3(new_n229), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n227), .A2(new_n245), .A3(new_n251), .A4(new_n229), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT82), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n248), .A2(new_n253), .A3(new_n260), .A4(new_n257), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n227), .A2(new_n229), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n246), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n255), .B1(new_n264), .B2(new_n249), .ZN(new_n265));
  INV_X1    g064(.A(new_n254), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n249), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n245), .B1(new_n227), .B2(new_n229), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n246), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n255), .B1(new_n273), .B2(new_n230), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n252), .A2(KEYINPUT78), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n250), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n249), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n259), .B(new_n261), .C1(new_n272), .C2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G85gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n276), .A2(new_n277), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n267), .B(new_n271), .C1(new_n288), .C2(new_n274), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n289), .A2(new_n284), .A3(new_n259), .A4(new_n261), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n279), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT22), .B1(new_n297), .B2(G218gat), .ZN(new_n298));
  XOR2_X1   g097(.A(G197gat), .B(G204gat), .Z(new_n299));
  OAI21_X1  g098(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G211gat), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n293), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(KEYINPUT27), .ZN(new_n311));
  AOI21_X1  g110(.A(G190gat), .B1(new_n310), .B2(KEYINPUT27), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(KEYINPUT27), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT28), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT67), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT28), .A4(new_n320), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n333), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n330), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(KEYINPUT23), .B2(new_n327), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n310), .A2(new_n320), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT65), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n327), .B2(KEYINPUT23), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n340), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n350), .A2(KEYINPUT64), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n350), .B2(KEYINPUT64), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n338), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n338), .B(KEYINPUT74), .C1(new_n352), .C2(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n308), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n358), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n360), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT64), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT25), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT64), .A3(new_n351), .ZN(new_n368));
  INV_X1    g167(.A(new_n337), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT68), .B1(new_n332), .B2(new_n333), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n367), .A2(new_n368), .B1(new_n371), .B2(new_n326), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n357), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n308), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n307), .A3(new_n373), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n361), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n308), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT37), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT38), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n385), .A3(new_n386), .A4(new_n377), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n291), .A2(new_n292), .A3(new_n379), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT90), .ZN(new_n389));
  INV_X1    g188(.A(new_n360), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n356), .B2(new_n358), .ZN(new_n391));
  INV_X1    g190(.A(new_n373), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n391), .A2(new_n392), .A3(new_n307), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n362), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n378), .B1(new_n394), .B2(new_n380), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT37), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n383), .B2(new_n308), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT38), .B1(new_n397), .B2(new_n382), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n395), .A2(new_n398), .B1(new_n394), .B2(new_n378), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n291), .A4(new_n292), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT37), .B1(new_n393), .B2(new_n362), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n386), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n300), .B2(new_n306), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n263), .B1(new_n412), .B2(KEYINPUT3), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n247), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n413), .A2(new_n414), .B1(new_n416), .B2(new_n308), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT84), .B(new_n263), .C1(new_n412), .C2(KEYINPUT3), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n411), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n307), .B1(new_n416), .B2(KEYINPUT85), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n247), .A2(new_n422), .A3(new_n415), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT86), .B(G22gat), .C1(new_n419), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n414), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n308), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n410), .ZN(new_n429));
  INV_X1    g228(.A(G22gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n308), .A3(new_n423), .ZN(new_n432));
  INV_X1    g231(.A(new_n420), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n434), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT86), .B1(new_n437), .B2(G22gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n409), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n419), .B2(new_n424), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n429), .A2(new_n434), .A3(new_n440), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n442), .A2(new_n408), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n264), .A2(new_n249), .A3(new_n255), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(KEYINPUT88), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(KEYINPUT88), .B2(new_n448), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n255), .B1(new_n248), .B2(new_n253), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n285), .B1(new_n451), .B2(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT40), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n279), .B2(new_n285), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n377), .B1(new_n393), .B2(new_n362), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n379), .A2(new_n459), .A3(KEYINPUT30), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n394), .A2(new_n461), .A3(new_n378), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n446), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n405), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n286), .A2(new_n467), .A3(new_n287), .A4(new_n290), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n279), .B(new_n285), .C1(KEYINPUT83), .C2(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n446), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n338), .B(new_n245), .C1(new_n352), .C2(new_n353), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n367), .A2(new_n368), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT70), .A3(new_n245), .A4(new_n338), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n354), .A2(new_n246), .ZN(new_n477));
  NAND2_X1  g276(.A1(G227gat), .A2(G233gat), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT32), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(new_n477), .A3(new_n476), .ZN(new_n484));
  INV_X1    g283(.A(new_n478), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT33), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AOI221_X4 g291(.A(new_n483), .B1(KEYINPUT33), .B2(new_n490), .C1(new_n484), .C2(new_n485), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n482), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n485), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n486), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n486), .B1(new_n487), .B2(new_n491), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n481), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n481), .B1(new_n499), .B2(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n494), .B2(new_n501), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n471), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n468), .A2(new_n469), .B1(new_n462), .B2(new_n460), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n446), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n515));
  INV_X1    g314(.A(new_n501), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n503), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n291), .A2(new_n292), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT35), .B1(new_n460), .B2(new_n462), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n446), .A4(new_n519), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n466), .A2(new_n512), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G15gat), .B(G22gat), .Z(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT92), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G8gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n528), .A2(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(G8gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n539), .A2(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n535), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n547), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n529), .B(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n546), .A3(new_n544), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n550), .A3(new_n557), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n552), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  INV_X1    g365(.A(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT11), .B(G169gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(new_n565), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n559), .B(new_n562), .C1(new_n564), .C2(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n202), .B1(new_n521), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n403), .B1(new_n388), .B2(KEYINPUT90), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n464), .B1(new_n579), .B2(new_n401), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n502), .B2(new_n505), .ZN(new_n582));
  OAI22_X1  g381(.A1(new_n582), .A2(new_n510), .B1(new_n446), .B2(new_n513), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n428), .A2(new_n410), .B1(new_n432), .B2(new_n433), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n430), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n435), .A3(new_n425), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n444), .B1(new_n588), .B2(new_n409), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n502), .B2(new_n505), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n584), .B1(new_n590), .B2(new_n513), .ZN(new_n591));
  INV_X1    g390(.A(new_n520), .ZN(new_n592));
  OAI22_X1  g391(.A1(new_n580), .A2(new_n583), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT96), .A3(new_n576), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n578), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G64gat), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n598), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G71gat), .ZN(new_n604));
  INV_X1    g403(.A(G78gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT97), .A3(new_n602), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT97), .B1(new_n606), .B2(new_n602), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n598), .A2(new_n600), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n601), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n602), .A3(new_n606), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n596), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n602), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n607), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n619), .B2(new_n603), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT21), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n531), .B(new_n534), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  AND2_X1   g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n631), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n632), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G99gat), .B(G106gat), .Z(new_n640));
  NAND2_X1  g439(.A1(G85gat), .A2(G92gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(G85gat), .A3(G92gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n644), .A3(KEYINPUT7), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT8), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(G99gat), .B2(G106gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT101), .B(G92gat), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n645), .B(new_n648), .C1(G85gat), .C2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT7), .B1(new_n642), .B2(new_n644), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n640), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT101), .B(G92gat), .Z(new_n653));
  INV_X1    g452(.A(G85gat), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n640), .ZN(new_n656));
  INV_X1    g455(.A(new_n651), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .A4(new_n645), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n554), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n548), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n666), .A3(new_n663), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  XNOR2_X1  g471(.A(G134gat), .B(G162gat), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n672), .B1(new_n671), .B2(new_n675), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n668), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n667), .A3(new_n676), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n639), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n658), .A2(KEYINPUT105), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n613), .B1(new_n618), .B2(new_n607), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n603), .A2(new_n616), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT98), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n610), .A2(new_n596), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n662), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n621), .A2(new_n659), .A3(new_n686), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT10), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n662), .A2(new_n621), .A3(KEYINPUT10), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n685), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n699), .B(new_n685), .C1(new_n694), .C2(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n691), .A2(new_n662), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n659), .B1(new_n621), .B2(new_n686), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n685), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(G120gat), .B(G148gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(G176gat), .B(G204gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n697), .ZN(new_n712));
  INV_X1    g511(.A(new_n706), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n684), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n595), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n470), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n523), .ZN(G1324gat));
  AND2_X1   g518(.A1(new_n595), .A2(new_n716), .ZN(new_n720));
  INV_X1    g519(.A(new_n463), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G8gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT16), .B(G8gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  MUX2_X1   g525(.A(new_n724), .B(KEYINPUT42), .S(new_n726), .Z(G1325gat));
  NAND2_X1  g526(.A1(new_n507), .A2(new_n511), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n720), .A2(G15gat), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(G15gat), .B1(new_n720), .B2(new_n517), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1326gat));
  NAND3_X1  g531(.A1(new_n720), .A2(new_n430), .A3(new_n589), .ZN(new_n733));
  OAI21_X1  g532(.A(G22gat), .B1(new_n717), .B2(new_n446), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  INV_X1    g536(.A(new_n639), .ZN(new_n738));
  INV_X1    g537(.A(new_n715), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n683), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n578), .A2(new_n594), .A3(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(G29gat), .A3(new_n470), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT45), .Z(new_n744));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n521), .B2(new_n683), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n593), .A2(new_n746), .A3(new_n682), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n740), .A2(new_n577), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n751), .B2(new_n470), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n744), .A2(new_n752), .ZN(G1328gat));
  OAI21_X1  g552(.A(G36gat), .B1(new_n751), .B2(new_n463), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n595), .A2(new_n538), .A3(new_n721), .A4(new_n741), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(new_n517), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n742), .A2(G43gat), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n748), .A2(new_n729), .A3(new_n749), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G43gat), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n760), .B2(new_n762), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT109), .B2(new_n765), .ZN(G1330gat));
  NAND3_X1  g566(.A1(new_n595), .A2(KEYINPUT110), .A3(new_n741), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n446), .B1(new_n742), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(G50gat), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n589), .A2(G50gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n750), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1331gat));
  NOR3_X1   g574(.A1(new_n684), .A2(new_n576), .A3(new_n739), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n593), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n470), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n597), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n463), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  OAI21_X1  g584(.A(new_n604), .B1(new_n778), .B2(new_n759), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n729), .A2(G71gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n778), .A2(new_n446), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n605), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n639), .A2(new_n576), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n715), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n593), .A2(new_n746), .A3(new_n682), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n746), .B1(new_n593), .B2(new_n682), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n748), .A2(KEYINPUT112), .A3(new_n794), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n470), .A2(new_n654), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n593), .A2(new_n682), .ZN(new_n804));
  INV_X1    g603(.A(new_n792), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n593), .A2(new_n792), .A3(KEYINPUT51), .A4(new_n682), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n470), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n715), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n801), .A2(new_n802), .B1(new_n810), .B2(new_n654), .ZN(G1336gat));
  NOR3_X1   g610(.A1(new_n739), .A2(G92gat), .A3(new_n463), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT113), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n649), .B1(new_n797), .B2(new_n463), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n807), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n817), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n748), .B2(new_n794), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n798), .B(new_n793), .C1(new_n745), .C2(new_n747), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n721), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n823), .B2(new_n649), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n817), .A2(new_n813), .A3(new_n819), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n463), .B1(new_n799), .B2(new_n800), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n653), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(KEYINPUT52), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n816), .B1(new_n826), .B2(new_n831), .ZN(G1337gat));
  NOR2_X1   g631(.A1(new_n759), .A2(G99gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n808), .A2(new_n715), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n801), .A2(KEYINPUT116), .A3(new_n729), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G99gat), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT116), .B1(new_n801), .B2(new_n729), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(G1338gat));
  AOI21_X1  g637(.A(new_n446), .B1(new_n799), .B2(new_n800), .ZN(new_n839));
  INV_X1    g638(.A(G106gat), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n589), .B1(new_n821), .B2(new_n822), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(G106gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n446), .A2(G106gat), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n817), .A2(new_n715), .A3(new_n819), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  OAI21_X1  g647(.A(G106gat), .B1(new_n797), .B2(new_n446), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n808), .A2(new_n715), .A3(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(G1339gat));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n710), .B1(new_n712), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n694), .A2(new_n696), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n856), .B2(new_n705), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT10), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n702), .B2(new_n703), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n695), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n699), .B1(new_n860), .B2(new_n685), .ZN(new_n861));
  INV_X1    g660(.A(new_n700), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT118), .B(new_n857), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT118), .B1(new_n701), .B2(new_n857), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT55), .B(new_n855), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(new_n576), .A3(new_n711), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n559), .A2(new_n562), .A3(new_n572), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n549), .A2(new_n551), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n570), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n715), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n682), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n868), .A2(new_n711), .A3(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n682), .A2(new_n875), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n738), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n639), .A2(new_n577), .A3(new_n683), .A4(new_n739), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n759), .A2(new_n589), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n470), .A2(new_n721), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G113gat), .B1(new_n889), .B2(new_n577), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n809), .A3(new_n590), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n721), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n235), .A3(new_n576), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(G1340gat));
  OAI21_X1  g693(.A(G120gat), .B1(new_n889), .B2(new_n739), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n236), .A3(new_n715), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1341gat));
  AOI21_X1  g696(.A(G127gat), .B1(new_n892), .B2(new_n639), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n738), .A2(new_n233), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n888), .B2(new_n899), .ZN(G1342gat));
  NAND2_X1  g699(.A1(new_n682), .A2(new_n463), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT119), .Z(new_n902));
  NOR3_X1   g701(.A1(new_n891), .A2(G134gat), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT56), .ZN(new_n904));
  OAI21_X1  g703(.A(G134gat), .B1(new_n889), .B2(new_n683), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1343gat));
  NAND2_X1  g705(.A1(new_n728), .A2(new_n886), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT120), .Z(new_n908));
  NAND2_X1  g707(.A1(new_n589), .A2(KEYINPUT57), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n877), .A2(KEYINPUT121), .B1(new_n878), .B2(new_n879), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n911), .B(new_n682), .C1(new_n870), .C2(new_n876), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n738), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n913), .B2(new_n882), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n446), .B1(new_n881), .B2(new_n882), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(KEYINPUT57), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n576), .B(new_n908), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT122), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n576), .A2(new_n205), .ZN(new_n920));
  NOR4_X1   g719(.A1(new_n919), .A2(new_n729), .A3(new_n887), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n917), .B2(G141gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n918), .A2(new_n922), .A3(KEYINPUT58), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT58), .ZN(new_n924));
  AOI221_X4 g723(.A(new_n921), .B1(KEYINPUT122), .B2(new_n924), .C1(new_n917), .C2(G141gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(G1344gat));
  OAI21_X1  g725(.A(new_n908), .B1(new_n914), .B2(new_n916), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(new_n739), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n206), .A2(new_n207), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(KEYINPUT59), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n933), .B(new_n446), .C1(new_n881), .C2(new_n882), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n739), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n908), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n937), .B2(G148gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n919), .A2(new_n729), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n886), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n715), .A2(new_n929), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n931), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1345gat));
  OR3_X1    g741(.A1(new_n927), .A2(new_n222), .A3(new_n738), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n222), .B1(new_n940), .B2(new_n738), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n927), .B2(new_n683), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n902), .A2(G162gat), .A3(new_n470), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1347gat));
  INV_X1    g748(.A(G169gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n885), .A2(new_n809), .A3(new_n463), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n576), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n590), .A2(new_n721), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n470), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n883), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(G169gat), .A3(new_n577), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n952), .A2(new_n958), .ZN(G1348gat));
  INV_X1    g758(.A(G176gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n739), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n883), .A2(new_n715), .A3(new_n956), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n951), .A2(new_n961), .B1(new_n960), .B2(new_n962), .ZN(G1349gat));
  INV_X1    g762(.A(new_n323), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n957), .A2(new_n964), .A3(new_n738), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n951), .A2(new_n639), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(G183gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT60), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n967), .B(new_n969), .ZN(G1350gat));
  AOI21_X1  g769(.A(new_n320), .B1(new_n951), .B2(new_n682), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT61), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n957), .A2(G190gat), .A3(new_n683), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n809), .A2(new_n463), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n728), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n919), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n567), .A3(new_n576), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n935), .A2(new_n976), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n567), .B1(new_n980), .B2(new_n576), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n979), .A2(new_n981), .ZN(G1352gat));
  INV_X1    g781(.A(new_n976), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n936), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  INV_X1    g784(.A(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n977), .A2(new_n986), .A3(new_n715), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT126), .B1(new_n987), .B2(KEYINPUT62), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n987), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n989));
  OAI221_X1 g788(.A(new_n985), .B1(KEYINPUT62), .B2(new_n987), .C1(new_n988), .C2(new_n989), .ZN(G1353gat));
  NAND3_X1  g789(.A1(new_n977), .A2(new_n302), .A3(new_n639), .ZN(new_n991));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n639), .B(new_n983), .C1(new_n916), .C2(new_n934), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(KEYINPUT127), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n916), .A2(new_n934), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n639), .A4(new_n983), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n994), .A2(new_n997), .A3(KEYINPUT63), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n994), .B2(new_n997), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(G1354gat));
  AOI21_X1  g799(.A(G218gat), .B1(new_n977), .B2(new_n682), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n683), .A2(new_n303), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n980), .B2(new_n1002), .ZN(G1355gat));
endmodule


