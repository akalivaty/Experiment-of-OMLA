//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n217), .B(new_n222), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(new_n205), .A2(G20), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT8), .A2(G58), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT8), .A2(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n220), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n257), .A2(new_n220), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G1), .B2(new_n212), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(G50), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n211), .C1(G41), .C2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n274), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G222), .A2(G1698), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT67), .B(G223), .Z(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G1698), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(G200), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n268), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(new_n251), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n211), .B2(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n261), .A2(new_n258), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n261), .B2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n252), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n212), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT7), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT7), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n306), .A3(new_n212), .A4(new_n303), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(G68), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(G58), .B(G68), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n263), .B1(new_n313), .B2(KEYINPUT16), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT74), .B1(new_n308), .B2(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n300), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n270), .A2(G232), .A3(new_n272), .A4(new_n274), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n320));
  INV_X1    g0120(.A(new_n220), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n269), .A2(KEYINPUT66), .B1(new_n321), .B2(new_n273), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(G232), .A4(new_n272), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G223), .B2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G87), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n327), .A2(new_n283), .B1(new_n252), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n274), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n279), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(G179), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT18), .B1(new_n318), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n258), .B1(new_n315), .B2(new_n316), .ZN(new_n337));
  AOI211_X1 g0137(.A(KEYINPUT74), .B(KEYINPUT16), .C1(new_n308), .C2(new_n310), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n299), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G169), .B1(new_n325), .B2(new_n331), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n325), .A2(new_n331), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  AOI21_X1  g0146(.A(G200), .B1(new_n325), .B2(new_n331), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n291), .B2(new_n342), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n346), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n314), .A2(new_n317), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n325), .A2(new_n291), .A3(new_n331), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n342), .B2(G200), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT17), .A4(new_n299), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n336), .A2(new_n345), .A3(new_n349), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  INV_X1    g0156(.A(new_n267), .ZN(new_n357));
  INV_X1    g0157(.A(new_n290), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n267), .B(KEYINPUT69), .C1(G169), .C2(new_n358), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(G179), .C2(new_n290), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n270), .A2(G244), .A3(new_n272), .A4(new_n274), .ZN(new_n363));
  INV_X1    g0163(.A(new_n279), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(G232), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n367));
  OAI211_X1 g0167(.A(G238), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n302), .A2(new_n303), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n208), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n330), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n291), .ZN(new_n373));
  OR2_X1    g0173(.A1(KEYINPUT8), .A2(G58), .ZN(new_n374));
  NAND2_X1  g0174(.A1(KEYINPUT8), .A2(G58), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n254), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n212), .A2(new_n284), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT70), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(new_n381), .A3(new_n378), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n253), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n258), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n260), .A2(G77), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n264), .B2(new_n284), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n365), .B2(new_n371), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n373), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n372), .A2(G179), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n390), .B1(new_n386), .B2(new_n258), .ZN(new_n397));
  AOI21_X1  g0197(.A(G169), .B1(new_n365), .B2(new_n371), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT71), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n395), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n295), .A2(new_n355), .A3(new_n362), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  OAI211_X1 g0205(.A(G226), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT72), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n369), .A2(new_n408), .A3(G226), .A4(new_n366), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n369), .A2(G232), .A3(G1698), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n330), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n275), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n322), .A2(KEYINPUT73), .A3(new_n272), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(G238), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n405), .A2(new_n413), .A3(new_n417), .A4(new_n364), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n279), .B1(new_n412), .B2(new_n330), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n405), .B1(new_n419), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g0220(.A(G200), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n417), .A3(new_n364), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n405), .A3(new_n417), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G190), .A3(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n426));
  INV_X1    g0226(.A(G50), .ZN(new_n427));
  INV_X1    g0227(.A(new_n254), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n429), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT11), .B1(new_n429), .B2(new_n258), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT12), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n261), .B2(new_n202), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n264), .A2(new_n202), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n430), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n421), .A2(new_n425), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n418), .B2(new_n420), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(G169), .C1(new_n418), .C2(new_n420), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n423), .A2(G179), .A3(new_n424), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n436), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n404), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n261), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n211), .A2(G33), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n263), .A2(new_n260), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(new_n449), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n257), .A2(new_n220), .B1(G20), .B2(new_n449), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(G33), .B2(G283), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n252), .A2(G97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT83), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT83), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(KEYINPUT20), .B(new_n454), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n453), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n211), .B(G45), .C1(new_n465), .C2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT77), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(KEYINPUT77), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n278), .B1(KEYINPUT5), .B2(new_n465), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n468), .A2(new_n473), .A3(new_n274), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G270), .A3(new_n274), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n302), .A2(G303), .A3(new_n303), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n330), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(G179), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n464), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n475), .A3(new_n478), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n453), .ZN(new_n490));
  INV_X1    g0290(.A(new_n463), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n455), .A2(new_n456), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n457), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n495), .B2(new_n454), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n490), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n479), .A2(KEYINPUT82), .A3(new_n484), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n489), .A2(new_n497), .A3(G169), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n486), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n487), .A2(new_n488), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT82), .B1(new_n479), .B2(new_n484), .ZN(new_n503));
  OAI21_X1  g0303(.A(G190), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n489), .A2(G200), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n464), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(KEYINPUT21), .A3(G169), .A4(new_n497), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n501), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n305), .A2(G107), .A3(new_n307), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT6), .A2(G97), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT76), .B1(new_n511), .B2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT76), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(new_n208), .A3(KEYINPUT6), .A4(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT6), .B1(new_n209), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(G20), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n254), .A2(G77), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n258), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n261), .A2(new_n207), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n452), .B2(new_n207), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT79), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n526), .B(new_n523), .C1(new_n520), .C2(new_n258), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n369), .A2(KEYINPUT4), .A3(G244), .A4(new_n366), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n369), .A2(G250), .A3(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n330), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n471), .A2(G41), .ZN(new_n536));
  OAI211_X1 g0336(.A(G257), .B(new_n274), .C1(new_n466), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n477), .A2(new_n539), .A3(G257), .A4(new_n274), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n474), .A2(new_n274), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT77), .B1(new_n470), .B2(new_n472), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n538), .A2(new_n540), .B1(new_n543), .B2(new_n473), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n535), .A2(new_n544), .A3(G179), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n333), .B1(new_n535), .B2(new_n544), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n525), .A2(new_n527), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n523), .B1(new_n520), .B2(new_n258), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n535), .A2(new_n544), .A3(G190), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n535), .A2(new_n544), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n393), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G116), .ZN(new_n552));
  OAI211_X1 g0352(.A(G238), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n330), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n211), .A2(G45), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n559), .A2(G250), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n274), .B1(new_n470), .B2(G274), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n333), .ZN(new_n563));
  INV_X1    g0363(.A(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n554), .A2(new_n555), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n369), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n552), .A4(new_n553), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n567), .B2(new_n330), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n341), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(new_n302), .B2(new_n303), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n253), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(G68), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n212), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n577), .A3(new_n212), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n328), .A2(new_n207), .A3(new_n208), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n263), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n452), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n384), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n384), .A2(new_n260), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n563), .A2(new_n569), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n452), .A2(new_n328), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n581), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n558), .A2(G190), .A3(new_n561), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n393), .C2(new_n568), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n547), .A2(new_n551), .A3(new_n588), .A4(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n212), .B(G87), .C1(new_n281), .C2(new_n282), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT22), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT22), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n369), .A2(new_n596), .A3(new_n212), .A4(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n552), .A2(G20), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n212), .B2(G107), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n599), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n258), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT25), .ZN(new_n609));
  AOI211_X1 g0409(.A(G107), .B(new_n260), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(G107), .B2(new_n583), .ZN(new_n614));
  OAI211_X1 g0414(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n615));
  OAI211_X1 g0415(.A(G250), .B(new_n366), .C1(new_n281), .C2(new_n282), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G294), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n330), .ZN(new_n619));
  OAI211_X1 g0419(.A(G264), .B(new_n274), .C1(new_n466), .C2(new_n536), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n475), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n477), .A2(KEYINPUT85), .A3(G264), .A4(new_n274), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n625), .B1(new_n618), .B2(new_n330), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(G179), .A3(new_n475), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n607), .A2(new_n614), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n607), .A2(new_n614), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n619), .A2(new_n621), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n625), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n618), .A2(new_n330), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n475), .A3(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n291), .A2(new_n631), .B1(new_n634), .B2(new_n393), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n629), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n393), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n633), .A2(new_n291), .A3(new_n475), .A4(new_n620), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(KEYINPUT86), .A3(new_n607), .A4(new_n614), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n628), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n448), .A2(new_n509), .A3(new_n593), .A4(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n588), .ZN(new_n643));
  INV_X1    g0443(.A(new_n547), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n588), .A2(new_n592), .ZN(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n588), .A2(new_n592), .ZN(new_n650));
  INV_X1    g0450(.A(new_n548), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n545), .B2(new_n546), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n643), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n636), .A2(new_n640), .ZN(new_n655));
  INV_X1    g0455(.A(new_n628), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n501), .A2(new_n656), .A3(new_n508), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n593), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n448), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n336), .A2(new_n345), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n437), .A2(new_n349), .A3(new_n353), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n333), .B1(new_n423), .B2(new_n424), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n443), .B1(new_n663), .B2(new_n441), .ZN(new_n664));
  INV_X1    g0464(.A(new_n442), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n445), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n401), .A2(new_n402), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n295), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n362), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n660), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n509), .B1(new_n464), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n501), .A2(new_n508), .ZN(new_n678));
  INV_X1    g0478(.A(new_n676), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n497), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT88), .Z(new_n682));
  NAND2_X1  g0482(.A1(new_n630), .A2(new_n679), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n641), .A2(new_n683), .B1(new_n628), .B2(new_n679), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(G330), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n641), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n679), .B1(new_n501), .B2(new_n508), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n676), .B(KEYINPUT89), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n656), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n215), .A2(new_n465), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n579), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n218), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n691), .B1(new_n654), .B2(new_n658), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n588), .B(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n652), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n645), .A2(KEYINPUT26), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n646), .B1(new_n650), .B2(new_n547), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n658), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n487), .A2(new_n341), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n550), .A2(new_n713), .A3(new_n568), .A4(new_n626), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n485), .A2(new_n562), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n550), .A4(new_n626), .ZN(new_n718));
  AOI21_X1  g0518(.A(G179), .B1(new_n535), .B2(new_n544), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n568), .B1(new_n475), .B2(new_n626), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n507), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n679), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n691), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n509), .A2(new_n593), .A3(new_n641), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n712), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n701), .B1(new_n732), .B2(G1), .ZN(G364));
  AND2_X1   g0533(.A1(new_n212), .A2(G13), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n211), .B1(new_n734), .B2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n697), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n682), .B2(G330), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G330), .B2(new_n682), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n215), .A2(new_n369), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n741), .B1(G116), .B2(new_n215), .ZN(new_n742));
  INV_X1    g0542(.A(new_n215), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n369), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n469), .B2(new_n219), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n243), .A2(new_n469), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n220), .B1(G20), .B2(new_n333), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n737), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n212), .B1(new_n756), .B2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n393), .A2(G179), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n212), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n369), .B1(new_n757), .B2(new_n207), .C1(new_n208), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n341), .A2(new_n393), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n341), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n202), .B1(new_n765), .B2(new_n284), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(new_n291), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n764), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n758), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n201), .A2(new_n768), .B1(new_n769), .B2(new_n328), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n761), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(new_n756), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT32), .ZN(new_n775));
  AND3_X1   g0575(.A1(new_n767), .A2(new_n762), .A3(KEYINPUT92), .ZN(new_n776));
  AOI21_X1  g0576(.A(KEYINPUT92), .B1(new_n767), .B2(new_n762), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n771), .B(new_n775), .C1(new_n427), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n283), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT93), .Z(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n760), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G317), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(KEYINPUT33), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(KEYINPUT33), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n763), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n768), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n784), .B(new_n788), .C1(G322), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G326), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  INV_X1    g0593(.A(G329), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n765), .A2(new_n793), .B1(new_n772), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n757), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(G294), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n790), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n779), .B1(new_n782), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n755), .B1(new_n799), .B2(new_n752), .ZN(new_n800));
  INV_X1    g0600(.A(new_n751), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n681), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n739), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  INV_X1    g0604(.A(new_n752), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n750), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n737), .B1(G77), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n283), .B1(new_n769), .B2(new_n208), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT95), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n791), .A2(G303), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n783), .A2(new_n763), .B1(new_n768), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n760), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G87), .B2(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n765), .A2(new_n449), .B1(new_n772), .B2(new_n793), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G97), .B2(new_n796), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n810), .A2(new_n811), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n765), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n789), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n763), .C1(new_n778), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n369), .B1(new_n769), .B2(new_n427), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n760), .A2(new_n202), .B1(new_n772), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(G58), .C2(new_n796), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n818), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n808), .B1(new_n752), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n372), .A2(new_n333), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n392), .A2(new_n834), .A3(new_n400), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n397), .A2(new_n676), .ZN(new_n836));
  INV_X1    g0636(.A(new_n396), .ZN(new_n837));
  AND4_X1   g0637(.A1(new_n402), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n403), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n833), .B1(new_n841), .B2(new_n750), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT96), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n702), .B(new_n840), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n730), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n730), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n844), .A2(KEYINPUT96), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(new_n736), .C1(new_n848), .C2(new_n844), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n847), .B2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT98), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n339), .A2(new_n675), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n354), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n350), .A2(new_n352), .A3(new_n299), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n339), .A2(new_n343), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n857), .A2(new_n858), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n354), .B2(new_n855), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n354), .A2(new_n855), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n852), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(KEYINPUT98), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n856), .A4(new_n863), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n852), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n444), .A2(new_n445), .A3(new_n676), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n436), .A2(new_n676), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n666), .A2(new_n437), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT97), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n446), .A2(KEYINPUT97), .A3(new_n881), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n884), .A2(new_n885), .B1(new_n444), .B2(new_n880), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n667), .A2(new_n679), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n702), .B2(new_n841), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n675), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n889), .A2(new_n874), .B1(new_n661), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n879), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n448), .A2(new_n703), .A3(new_n711), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n670), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n892), .B(new_n894), .Z(new_n895));
  INV_X1    g0695(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n863), .A2(new_n868), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n865), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n873), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n873), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n728), .A2(new_n726), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n841), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n886), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n444), .A2(new_n880), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n882), .A2(new_n883), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT97), .B1(new_n446), .B2(new_n881), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n904), .A2(new_n841), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n874), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n901), .A2(new_n906), .B1(new_n912), .B2(new_n902), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n448), .A2(new_n904), .ZN(new_n915));
  OAI21_X1  g0715(.A(G330), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n914), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n895), .A2(new_n917), .B1(new_n211), .B2(new_n734), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n895), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n515), .A2(new_n517), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(G116), .A3(new_n221), .A4(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  OAI211_X1 g0725(.A(new_n219), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n427), .A2(G68), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n211), .B(G13), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n919), .A2(new_n925), .A3(new_n928), .ZN(G367));
  NOR2_X1   g0729(.A1(new_n769), .A2(new_n449), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n369), .B(new_n931), .C1(G303), .C2(new_n789), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n930), .A2(KEYINPUT46), .B1(G107), .B2(new_n796), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n791), .A2(G311), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n207), .A2(new_n760), .B1(new_n765), .B2(new_n783), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n763), .A2(new_n812), .B1(new_n772), .B2(new_n785), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n763), .A2(new_n773), .B1(new_n772), .B2(new_n822), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n369), .B1(new_n769), .B2(new_n201), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n757), .A2(new_n202), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(G150), .A2(new_n789), .B1(new_n819), .B2(G50), .ZN(new_n943));
  INV_X1    g0743(.A(G143), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n284), .B2(new_n760), .C1(new_n778), .C2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n938), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT105), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n752), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n590), .A2(new_n676), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n650), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n643), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n751), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n744), .A2(new_n239), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n754), .B1(new_n743), .B2(new_n384), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n736), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n690), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n547), .B(new_n551), .C1(new_n548), .C2(new_n727), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n706), .A2(new_n691), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n958), .A2(KEYINPUT42), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n547), .B1(new_n962), .B2(new_n656), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n727), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT42), .B1(new_n958), .B2(new_n962), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT100), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT100), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n951), .A2(new_n952), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT43), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT101), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(KEYINPUT101), .A3(new_n972), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n968), .A2(new_n969), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n686), .A2(new_n962), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n735), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n961), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT104), .B1(new_n693), .B2(new_n961), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n693), .A2(new_n961), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n686), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n682), .A2(G330), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n690), .B1(new_n684), .B2(new_n689), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n988), .A2(new_n686), .A3(new_n989), .A4(new_n992), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n732), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n732), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n697), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n983), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n957), .B1(new_n982), .B2(new_n1004), .ZN(G387));
  OR2_X1    g0805(.A1(new_n998), .A2(new_n732), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n998), .A2(new_n732), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n697), .B(KEYINPUT110), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n684), .A2(new_n751), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n740), .A2(new_n698), .B1(G107), .B2(new_n215), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n745), .B1(new_n236), .B2(G45), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n698), .B(new_n469), .C1(new_n202), .C2(new_n284), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n296), .B2(G50), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n296), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1011), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n737), .B1(new_n1019), .B2(new_n754), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n769), .A2(new_n284), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G68), .B2(new_n819), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n821), .B2(new_n772), .C1(new_n296), .C2(new_n763), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n283), .B(new_n1023), .C1(G97), .C2(new_n814), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n757), .A2(new_n383), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G50), .B2(new_n789), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT107), .Z(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n1027), .C1(new_n773), .C2(new_n778), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT108), .Z(new_n1029));
  INV_X1    g0829(.A(new_n772), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n369), .B1(new_n1030), .B2(G326), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n789), .B1(new_n819), .B2(G303), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n763), .A2(new_n793), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n791), .B2(G322), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1035), .A2(KEYINPUT109), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(KEYINPUT109), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n769), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1042), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1031), .B1(new_n449), .B2(new_n760), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1029), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1020), .B1(new_n1048), .B2(new_n752), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n998), .A2(new_n983), .B1(new_n1010), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1009), .A2(new_n1050), .ZN(G393));
  INV_X1    g0851(.A(KEYINPUT111), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n995), .B2(new_n999), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n999), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1007), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1000), .B(new_n1008), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n962), .A2(new_n751), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n753), .B1(new_n207), .B2(new_n215), .C1(new_n745), .C2(new_n246), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n737), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n778), .A2(new_n821), .B1(new_n773), .B2(new_n768), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT113), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G68), .A2(new_n1042), .B1(new_n1030), .B2(G143), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n427), .B2(new_n763), .C1(new_n296), .C2(new_n765), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n796), .A2(G77), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n369), .C1(new_n328), .C2(new_n760), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n785), .B1(new_n793), .B2(new_n768), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  AOI22_X1  g0870(.A1(G283), .A2(new_n1042), .B1(new_n1030), .B2(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n812), .B2(new_n765), .C1(new_n780), .C2(new_n763), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n283), .B1(new_n757), .B2(new_n449), .C1(new_n208), .C2(new_n760), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1059), .B1(new_n1075), .B2(new_n752), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1054), .A2(new_n983), .B1(new_n1057), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1056), .A2(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(KEYINPUT114), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n679), .B(new_n840), .C1(new_n709), .C2(new_n658), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n887), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n710), .A2(new_n676), .A3(new_n841), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n887), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(KEYINPUT114), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n910), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT99), .B1(new_n867), .B2(new_n869), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n873), .A2(new_n898), .A3(new_n896), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1085), .A2(new_n877), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n877), .B1(new_n886), .B2(new_n888), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n874), .A2(new_n852), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT39), .B1(new_n873), .B2(new_n898), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n848), .A2(new_n910), .A3(new_n841), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n884), .A2(new_n885), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n905), .B1(new_n1095), .B2(new_n907), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(G330), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n910), .A2(G330), .A3(new_n911), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1088), .A2(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n875), .A2(new_n749), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n737), .B1(new_n251), .B2(new_n806), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT116), .Z(new_n1105));
  OAI22_X1  g0905(.A1(new_n202), .A2(new_n760), .B1(new_n765), .B2(new_n207), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n369), .B(new_n1106), .C1(G87), .C2(new_n1042), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n791), .A2(G283), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n208), .A2(new_n763), .B1(new_n768), .B2(new_n449), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G294), .B2(new_n1030), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1066), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n791), .A2(G128), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n769), .A2(new_n821), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n369), .B1(new_n760), .B2(new_n427), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G159), .B2(new_n796), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n827), .A2(new_n768), .B1(new_n763), .B2(new_n822), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n765), .A2(new_n1118), .B1(new_n772), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .A4(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1111), .A2(KEYINPUT117), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT117), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n805), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1105), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1102), .A2(new_n983), .B1(new_n1103), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n448), .A2(G330), .A3(new_n904), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n893), .A2(new_n1128), .A3(new_n670), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n886), .B1(new_n730), .B2(new_n840), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1100), .A2(new_n1098), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n888), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n904), .A2(G330), .A3(new_n841), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n886), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1134), .A2(new_n1093), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1129), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1008), .B1(new_n1102), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n899), .A2(new_n900), .A3(new_n878), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1142), .A2(new_n1085), .B1(new_n875), .B2(new_n1089), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1100), .A2(new_n1098), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1137), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1145), .A2(new_n1129), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1127), .B1(new_n1140), .B2(new_n1147), .ZN(G378));
  INV_X1    g0948(.A(KEYINPUT120), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n879), .B2(new_n891), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n357), .A2(new_n890), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n295), .B2(new_n362), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n295), .A2(new_n362), .A3(new_n1153), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n913), .B2(G330), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n912), .A2(new_n902), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1086), .A2(new_n1096), .A3(KEYINPUT40), .A4(new_n1087), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1161), .A4(G330), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1160), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1164), .A3(G330), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1168), .B2(KEYINPUT119), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1151), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(KEYINPUT119), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n1165), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1174), .A2(new_n1150), .A3(new_n1169), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n983), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n737), .B1(G50), .B2(new_n806), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n763), .A2(new_n827), .B1(new_n765), .B2(new_n822), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1179), .A2(new_n768), .B1(new_n769), .B2(new_n1118), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G150), .C2(new_n796), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1119), .B2(new_n778), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n814), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n1030), .C2(G124), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G50), .B1(new_n303), .B2(new_n465), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n814), .A2(G58), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT118), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n207), .A2(new_n763), .B1(new_n768), .B2(new_n208), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n765), .A2(new_n383), .B1(new_n772), .B2(new_n783), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n791), .A2(G116), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1021), .A2(new_n941), .A3(G41), .A4(new_n369), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1190), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1188), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1187), .B(new_n1198), .C1(new_n1197), .C2(new_n1196), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1177), .B1(new_n1199), .B2(new_n752), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1172), .B2(new_n750), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1129), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT57), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1174), .A2(new_n892), .A3(new_n1169), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT121), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n892), .B1(new_n1174), .B2(new_n1169), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT121), .B(new_n892), .C1(new_n1174), .C2(new_n1169), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1129), .B1(new_n1102), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1167), .A2(new_n1170), .A3(new_n1151), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1150), .B1(new_n1174), .B2(new_n1169), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1008), .B1(new_n1215), .B2(KEYINPUT57), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1176), .B(new_n1201), .C1(new_n1210), .C2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1211), .A2(new_n1202), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1133), .A2(new_n1129), .A3(new_n1138), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1003), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT122), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1190), .B1(new_n827), .B2(new_n778), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n757), .A2(new_n427), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n369), .B1(new_n768), .B2(new_n822), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n763), .A2(new_n1118), .B1(new_n765), .B2(new_n821), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n769), .A2(new_n773), .B1(new_n772), .B2(new_n1179), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT123), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n763), .A2(new_n449), .B1(new_n772), .B2(new_n780), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n283), .B1(new_n760), .B2(new_n284), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1025), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G97), .A2(new_n1042), .B1(new_n789), .B2(G283), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n208), .B2(new_n765), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n791), .B2(G294), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1226), .A2(new_n1228), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n737), .B1(G68), .B2(new_n806), .C1(new_n1235), .C2(new_n805), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n886), .B2(new_n749), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1211), .B2(new_n983), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1221), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G381));
  NAND3_X1  g1040(.A1(new_n1009), .A2(new_n803), .A3(new_n1050), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G384), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1056), .A3(new_n1077), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G387), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1239), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G407));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT125), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(new_n1251), .C2(new_n1254), .ZN(G409));
  OAI211_X1 g1055(.A(new_n1127), .B(new_n1201), .C1(new_n1140), .C2(new_n1147), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1003), .B2(new_n1215), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1207), .A2(new_n1206), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1167), .A2(new_n879), .A3(new_n891), .A4(new_n1170), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1209), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n983), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1250), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1176), .A2(new_n1201), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1008), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1203), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT57), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1204), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1263), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1262), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1250), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1219), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1129), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1218), .A3(new_n1008), .A4(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(new_n1238), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1277), .B2(new_n1238), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1273), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1238), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1277), .A2(G384), .A3(new_n1238), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1273), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G375), .A2(G378), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .A4(new_n1262), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1262), .B(new_n1291), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1288), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G393), .A2(G396), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n1241), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1241), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1056), .A3(new_n1077), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(G387), .ZN(new_n1302));
  INV_X1    g1102(.A(G387), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1295), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(KEYINPUT61), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1289), .A2(KEYINPUT63), .A3(new_n1291), .A4(new_n1262), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1280), .A2(new_n1286), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1309), .B1(new_n1313), .B2(new_n1272), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1293), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1307), .B(new_n1308), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1306), .A2(new_n1316), .ZN(G405));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1289), .A2(new_n1319), .A3(new_n1291), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1291), .B1(new_n1289), .B2(new_n1319), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1318), .B(new_n1305), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1322), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1305), .A2(new_n1318), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1302), .A2(KEYINPUT127), .A3(new_n1304), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1320), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1323), .A2(new_n1327), .ZN(G402));
endmodule


