//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G137), .A4(new_n465), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n462), .A2(new_n464), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND4_X1   g066(.A1(G126), .A2(new_n462), .A3(new_n464), .A4(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT69), .A2(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n497), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(KEYINPUT70), .C1(new_n495), .C2(new_n494), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n492), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(new_n504), .A3(G138), .A4(new_n465), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n513), .A2(new_n515), .A3(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(G651), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n522), .B1(new_n519), .B2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(G88), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(new_n522), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(new_n537), .A3(new_n525), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(G543), .A3(new_n537), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n523), .A2(KEYINPUT73), .A3(G543), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n539), .B1(G51), .B2(new_n544), .ZN(G168));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n538), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n513), .A2(new_n515), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n548), .A2(G90), .B1(G651), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n547), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n538), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n544), .B2(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n550), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n548), .A2(G91), .B1(G651), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT75), .B(KEYINPUT9), .Z(new_n573));
  NAND4_X1  g148(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n540), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n527), .B(new_n580), .ZN(G303));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n523), .A2(KEYINPUT77), .A3(G49), .A4(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n523), .A2(G87), .A3(new_n525), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n550), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n523), .A2(G48), .A3(G543), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n538), .ZN(G305));
  XNOR2_X1  g170(.A(KEYINPUT78), .B(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n548), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n542), .A2(new_n543), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI221_X1 g175(.A(new_n597), .B1(new_n521), .B2(new_n598), .C1(new_n599), .C2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G171), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n538), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .A4(new_n525), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n521), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n542), .A2(G54), .A3(new_n543), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n609), .A2(new_n612), .A3(KEYINPUT80), .A4(new_n611), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(KEYINPUT79), .B2(new_n603), .ZN(G284));
  OAI21_X1  g195(.A(new_n619), .B1(KEYINPUT79), .B2(new_n603), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n602), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n617), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n617), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n468), .A2(new_n478), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT13), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n484), .A2(G123), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT83), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n486), .A2(G135), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT82), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n640), .A2(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(new_n640), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n635), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G2438), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n651), .B(new_n652), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n665), .B2(new_n666), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n677), .A2(KEYINPUT17), .A3(new_n674), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n677), .B2(KEYINPUT17), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n678), .A2(new_n679), .A3(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n684), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n686), .A2(new_n684), .A3(new_n689), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n692), .A3(new_n689), .ZN(new_n694));
  AND4_X1   g269(.A1(new_n690), .A2(new_n691), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1991), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n697), .A2(G1996), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(G1996), .B1(new_n697), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n700), .B2(new_n701), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n705), .ZN(new_n708));
  INV_X1    g283(.A(new_n702), .ZN(new_n709));
  INV_X1    g284(.A(new_n701), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n708), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n712), .ZN(G229));
  NAND2_X1  g288(.A1(G288), .A2(KEYINPUT92), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n587), .A2(new_n586), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n715), .A2(new_n716), .A3(new_n585), .A4(new_n584), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G23), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n719), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G6), .B(G305), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n724), .A2(new_n725), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI22_X1  g311(.A1(G119), .A2(new_n484), .B1(new_n486), .B2(G131), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n738), .A2(G95), .A3(G2105), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(G95), .B2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n737), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G25), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT35), .B(G1991), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT90), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n743), .B(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n719), .A2(G24), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G290), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1986), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n746), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n735), .A2(new_n736), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n754));
  XOR2_X1   g329(.A(new_n753), .B(new_n754), .Z(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n483), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2105), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT97), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n478), .A2(G103), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT25), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT25), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n763), .A2(new_n764), .B1(G139), .B2(new_n486), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G33), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(G29), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n767), .B(new_n772), .C1(G29), .C2(new_n768), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT99), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT99), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n770), .A2(new_n773), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G2072), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n478), .A2(G105), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n484), .A2(G129), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n486), .A2(G141), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  AND4_X1   g361(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n781), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT27), .B(G1996), .Z(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT24), .ZN(new_n791));
  INV_X1    g366(.A(G34), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n481), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(G2084), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n780), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n777), .A2(new_n778), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n719), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n617), .B2(new_n719), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(G301), .A2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G5), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n814));
  INV_X1    g389(.A(G29), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n484), .A2(G128), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n486), .A2(G140), .ZN(new_n819));
  OR2_X1    g394(.A1(G104), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n824), .A2(KEYINPUT95), .A3(new_n815), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n822), .B(KEYINPUT94), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G29), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G2067), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n815), .A2(G27), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G164), .B2(new_n815), .ZN(new_n833));
  INV_X1    g408(.A(G2078), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G2084), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n788), .A2(new_n789), .B1(new_n796), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n815), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n815), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT29), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n835), .B(new_n837), .C1(G2090), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n719), .A2(G19), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n562), .B2(new_n719), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1341), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g420(.A1(new_n805), .A2(new_n813), .A3(new_n831), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n801), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n719), .A2(G20), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT23), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT23), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G299), .B2(G16), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n851), .B2(new_n848), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(G1956), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(G1956), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n840), .A2(G2090), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n777), .A2(new_n800), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(KEYINPUT100), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT30), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(G28), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n815), .B1(new_n863), .B2(G28), .ZN(new_n865));
  AND2_X1   g440(.A1(KEYINPUT31), .A2(G11), .ZN(new_n866));
  NOR2_X1   g441(.A1(KEYINPUT31), .A2(G11), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n864), .A2(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT85), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n645), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(new_n815), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n646), .A2(KEYINPUT102), .A3(G29), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n809), .A2(G1961), .A3(new_n810), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n719), .A2(G21), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G168), .B2(new_n719), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT101), .B(G1966), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT104), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n847), .A2(new_n862), .A3(KEYINPUT106), .A4(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n846), .A3(new_n801), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n799), .B1(new_n776), .B2(new_n775), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n859), .B(new_n858), .C1(new_n888), .C2(new_n778), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n755), .B1(new_n885), .B2(new_n890), .ZN(G311));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n885), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n753), .B(new_n754), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(G150));
  INV_X1    g469(.A(G93), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n538), .A2(new_n895), .B1(new_n896), .B2(new_n521), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n544), .B2(G55), .ZN(new_n898));
  INV_X1    g473(.A(G860), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n617), .A2(G559), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT39), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT107), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT38), .ZN(new_n905));
  INV_X1    g480(.A(G43), .ZN(new_n906));
  OAI221_X1 g481(.A(new_n559), .B1(new_n560), .B2(new_n538), .C1(new_n599), .C2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n898), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n899), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(G145));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n766), .B(new_n787), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n742), .B(new_n633), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n484), .A2(G130), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n486), .A2(G142), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n465), .A2(G118), .ZN(new_n918));
  OAI21_X1  g493(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n824), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n824), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G164), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n507), .A3(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n915), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n913), .A2(new_n914), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n913), .A2(new_n914), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n924), .A3(new_n925), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n871), .A2(G162), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n646), .A2(new_n490), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(G160), .ZN(new_n934));
  AOI21_X1  g509(.A(G160), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n912), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n935), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n933), .A3(G160), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(KEYINPUT108), .A3(new_n930), .A4(new_n927), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n931), .B2(new_n936), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g520(.A(new_n627), .B(new_n908), .ZN(new_n946));
  INV_X1    g521(.A(G299), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n613), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n613), .A2(G299), .A3(KEYINPUT109), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n952), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n946), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(G305), .B(new_n527), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n718), .B(G290), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n965), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n962), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n954), .A2(new_n960), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n963), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n963), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G868), .B2(new_n898), .ZN(G295));
  OAI21_X1  g553(.A(new_n977), .B1(G868), .B2(new_n898), .ZN(G331));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n967), .A2(new_n968), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n964), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n970), .ZN(new_n985));
  XNOR2_X1  g560(.A(G301), .B(G168), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(new_n908), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n908), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n959), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n956), .A3(new_n988), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(G37), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n984), .A2(new_n990), .A3(new_n970), .A4(new_n991), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n982), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n955), .A2(new_n958), .B1(new_n987), .B2(new_n988), .ZN(new_n997));
  INV_X1    g572(.A(new_n991), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n969), .A2(new_n971), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AND4_X1   g574(.A1(new_n996), .A2(new_n994), .A3(new_n999), .A4(new_n982), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n980), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n993), .A2(new_n982), .A3(new_n994), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n999), .A3(new_n996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(G397));
  AOI21_X1  g581(.A(G1384), .B1(new_n501), .B2(new_n506), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n472), .A2(new_n480), .A3(G40), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT45), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT114), .Z(new_n1010));
  INV_X1    g585(.A(new_n787), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n827), .A2(G2067), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n824), .A2(new_n830), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT46), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  OAI221_X1 g596(.A(new_n1016), .B1(new_n1011), .B2(new_n1018), .C1(new_n1012), .C2(new_n1017), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n742), .A2(new_n745), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n742), .A2(new_n745), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1010), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1009), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1021), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1024), .B(KEYINPUT125), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1014), .B1(new_n1022), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1010), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  INV_X1    g612(.A(G40), .ZN(new_n1038));
  NOR4_X1   g613(.A1(new_n471), .A2(new_n477), .A3(new_n1038), .A4(new_n479), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1041), .B(G1384), .C1(new_n501), .C2(new_n506), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(new_n1037), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1039), .B1(new_n1007), .B2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT50), .B(G1384), .C1(new_n501), .C2(new_n506), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n836), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1046), .A3(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1036), .B(G8), .C1(new_n1052), .C2(G286), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G168), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1036), .B(new_n1055), .C1(new_n1052), .C2(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT62), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(G8), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(KEYINPUT51), .C1(new_n1054), .C2(G168), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1056), .A4(new_n1053), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1054), .B1(new_n1039), .B2(new_n1007), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1064), .B(new_n1066), .C1(new_n718), .C2(new_n1065), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n714), .B2(new_n717), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1064), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G305), .A2(G1981), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n548), .A2(G86), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n593), .A4(new_n592), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1074), .A3(KEYINPUT49), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1064), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1067), .A2(new_n1070), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1384), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n507), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1008), .B1(new_n1082), .B2(new_n1041), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1007), .A2(KEYINPUT115), .A3(KEYINPUT45), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n728), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1050), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1054), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G303), .A2(G8), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1080), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1096), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1088), .A2(new_n728), .B1(new_n1050), .B2(new_n1090), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1054), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1083), .A2(new_n834), .A3(new_n1085), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1083), .A2(KEYINPUT123), .A3(new_n834), .A4(new_n1085), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT53), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1083), .A2(new_n1087), .A3(new_n834), .A4(new_n1084), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1049), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1082), .A2(KEYINPUT50), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n1039), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1109), .A2(new_n1110), .B1(new_n1113), .B2(new_n812), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1098), .A2(new_n1103), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1059), .A2(new_n1063), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n615), .A2(new_n616), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n804), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1039), .A2(new_n1007), .A3(new_n830), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1083), .A2(new_n1087), .A3(new_n1084), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT121), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G299), .B(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1121), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1124), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1119), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n1139), .B2(new_n1121), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n617), .A2(new_n1119), .A3(new_n1141), .A4(new_n1120), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT122), .B(G1996), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1083), .A2(new_n1087), .A3(new_n1084), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1039), .A2(new_n1007), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1143), .B1(new_n1149), .B2(new_n562), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT59), .B(new_n907), .C1(new_n1145), .C2(new_n1148), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1140), .B(new_n1142), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1135), .A2(KEYINPUT61), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1137), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1138), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(G301), .B(KEYINPUT54), .Z(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1050), .A2(KEYINPUT124), .A3(G1961), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT124), .B1(new_n1050), .B2(G1961), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT115), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1040), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1971), .B1(new_n1168), .B2(new_n1084), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1113), .A2(G2090), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1097), .B(G8), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1080), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1103), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1166), .B(new_n1174), .C1(new_n1058), .C2(new_n1057), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1117), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1052), .A2(G8), .A3(G168), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1178), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1098), .A2(new_n1180), .A3(KEYINPUT63), .A4(new_n1103), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(G288), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1079), .A2(new_n1065), .A3(new_n1183), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1184), .A2(new_n1074), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1185), .A2(new_n1069), .B1(new_n1171), .B2(new_n1080), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT117), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1189), .B(new_n1186), .C1(new_n1179), .C2(new_n1181), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1176), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  AND2_X1   g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT113), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1192), .A2(new_n1028), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(G290), .A2(new_n1193), .A3(G1986), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1009), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1023), .B(new_n1026), .C1(new_n1194), .C2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1035), .B1(new_n1191), .B2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g773(.A(new_n459), .B(G227), .C1(new_n667), .C2(new_n669), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n707), .A3(new_n712), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(KEYINPUT127), .ZN(new_n1202));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1203));
  NAND4_X1  g777(.A1(new_n1200), .A2(new_n1203), .A3(new_n707), .A4(new_n712), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n1202), .A2(new_n944), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1003), .A2(new_n981), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1206), .B2(new_n1002), .ZN(G308));
  NAND2_X1  g781(.A1(new_n1002), .A2(new_n1206), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n1208), .A2(new_n944), .A3(new_n1204), .A4(new_n1202), .ZN(G225));
endmodule


