//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n629, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT64), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(KEYINPUT65), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n462), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n459), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n470), .A2(new_n471), .A3(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT66), .B1(new_n459), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G101), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n475), .A2(G136), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT67), .Z(new_n481));
  NAND2_X1  g056(.A1(new_n460), .A2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n459), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n481), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT68), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n459), .C1(new_n464), .C2(new_n465), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n462), .A2(new_n466), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(KEYINPUT6), .B2(new_n506), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n506), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT69), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n509), .B(G651), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n503), .B1(new_n512), .B2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n507), .A2(new_n519), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n515), .B2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(KEYINPUT69), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n527), .B2(G651), .ZN(new_n528));
  AOI211_X1 g103(.A(KEYINPUT70), .B(new_n506), .C1(new_n525), .C2(new_n526), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT7), .Z(new_n538));
  AND3_X1   g113(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n539));
  AOI211_X1 g114(.A(new_n538), .B(new_n539), .C1(G89), .C2(new_n520), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n534), .A2(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n503), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(G90), .B1(G651), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n532), .B2(new_n533), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n503), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n520), .A2(G81), .B1(G651), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n503), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n512), .A2(new_n517), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  OAI211_X1 g146(.A(G53), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n518), .A2(new_n575), .A3(G53), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n573), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT74), .ZN(new_n580));
  AND4_X1   g155(.A1(new_n575), .A2(new_n567), .A3(G53), .A4(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n575), .B1(new_n518), .B2(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT73), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n570), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n580), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n506), .B1(new_n503), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n520), .B2(G87), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  AND2_X1   g167(.A1(G49), .A2(G543), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n567), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n592), .B1(new_n567), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(new_n520), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n518), .A2(G48), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n503), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n534), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n503), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n520), .A2(G85), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n520), .A2(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n532), .B2(new_n533), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n506), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n613), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n619));
  AOI211_X1 g194(.A(new_n531), .B(new_n508), .C1(new_n512), .C2(new_n517), .ZN(new_n620));
  OAI21_X1  g195(.A(G54), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n617), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(KEYINPUT76), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n612), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n610), .B1(new_n624), .B2(G868), .ZN(G321));
  MUX2_X1   g201(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g202(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n624), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g208(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  OR2_X1    g210(.A1(new_n472), .A2(new_n473), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n636), .A2(new_n466), .A3(new_n462), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n475), .A2(G135), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n459), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  INV_X1    g222(.A(G123), .ZN(new_n648));
  OAI221_X1 g223(.A(new_n645), .B1(new_n646), .B2(new_n647), .C1(new_n648), .C2(new_n483), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT80), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n642), .A2(new_n643), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2443), .B(G2446), .Z(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(G14), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n664), .ZN(G401));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n677), .B2(new_n671), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n671), .B(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n677), .A3(new_n674), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n676), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n687), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT83), .Z(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G171), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G5), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G1961), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  NAND2_X1  g284(.A1(G286), .A2(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G21), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT97), .B(G1966), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT99), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G33), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n475), .A2(G139), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n462), .A2(new_n466), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n722), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n459), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n716), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  OAI211_X1 g302(.A(new_n709), .B(new_n715), .C1(G2072), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n730), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n706), .A2(new_n707), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT85), .B(G16), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n557), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G19), .B2(new_n736), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n734), .B(new_n735), .C1(G1341), .C2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR2_X1   g316(.A1(new_n650), .A2(new_n716), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n741), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT24), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n716), .B1(new_n748), .B2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G160), .B2(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G2084), .ZN(new_n752));
  NOR2_X1   g327(.A1(G164), .A2(new_n716), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G27), .B2(new_n716), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2078), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n747), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n484), .A2(G129), .B1(new_n475), .B2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n636), .A2(G105), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT95), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n716), .B2(G32), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT27), .B(G1996), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n766), .A2(new_n768), .B1(G2078), .B2(new_n755), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n768), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n716), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G128), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n475), .A2(G140), .ZN(new_n775));
  OR2_X1    g350(.A1(G104), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(new_n716), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n770), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n751), .A2(G2084), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n757), .A2(new_n769), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n739), .A2(G1341), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(new_n712), .C2(new_n713), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n728), .A2(new_n740), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n727), .A2(G2072), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n704), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n624), .B2(new_n704), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n736), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1956), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n788), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n704), .A2(G23), .ZN(new_n807));
  INV_X1    g382(.A(G288), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n704), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(new_n805), .ZN(new_n812));
  INV_X1    g387(.A(new_n736), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(G22), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G166), .B2(new_n813), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT88), .B(G1971), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n806), .A2(new_n811), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n716), .A2(G25), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(G107), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G2105), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT84), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n475), .A2(G131), .ZN(new_n826));
  INV_X1    g401(.A(G119), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n483), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n821), .B1(new_n829), .B2(new_n716), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n813), .A2(G24), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G290), .B2(new_n736), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT86), .B(G1986), .Z(new_n835));
  OAI21_X1  g410(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n819), .A2(new_n820), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT89), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT89), .B(KEYINPUT36), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n801), .A2(new_n841), .A3(new_n844), .ZN(G311));
  INV_X1    g420(.A(G311), .ZN(G150));
  INV_X1    g421(.A(new_n612), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n615), .A2(new_n613), .A3(new_n617), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT76), .B1(new_n621), .B2(new_n622), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n629), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  OAI21_X1  g427(.A(G43), .B1(new_n619), .B2(new_n620), .ZN(new_n853));
  OAI21_X1  g428(.A(G55), .B1(new_n619), .B2(new_n620), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n503), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n520), .A2(G93), .B1(G651), .B2(new_n857), .ZN(new_n858));
  AND4_X1   g433(.A1(new_n853), .A2(new_n854), .A3(new_n555), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n853), .A2(new_n555), .B1(new_n854), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n852), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n532), .B2(new_n533), .ZN(new_n867));
  INV_X1    g442(.A(new_n858), .ZN(new_n868));
  OAI21_X1  g443(.A(G860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(new_n725), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n494), .A2(KEYINPUT103), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n490), .A2(new_n493), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n873), .A2(new_n875), .B1(new_n496), .B2(new_n499), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n778), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n764), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n764), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n641), .A2(new_n829), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n829), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n484), .A2(G130), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n475), .A2(G142), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT104), .ZN(new_n890));
  OR2_X1    g465(.A1(G106), .A2(G2105), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n891), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n885), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n885), .B2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n882), .A2(new_n898), .A3(KEYINPUT106), .A4(new_n883), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n882), .A2(new_n883), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n897), .B(new_n899), .C1(KEYINPUT106), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n650), .B(G160), .ZN(new_n902));
  XOR2_X1   g477(.A(G162), .B(new_n902), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n896), .A2(KEYINPUT107), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n882), .A2(new_n883), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n882), .B2(new_n883), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(new_n903), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n905), .A2(new_n913), .A3(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT40), .B1(new_n905), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(G395));
  XNOR2_X1  g491(.A(G290), .B(G303), .ZN(new_n917));
  XOR2_X1   g492(.A(G288), .B(G305), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n920), .B2(KEYINPUT110), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(KEYINPUT42), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(KEYINPUT42), .B2(new_n921), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n631), .B(new_n861), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n583), .A2(new_n584), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n586), .B1(new_n927), .B2(new_n571), .ZN(new_n928));
  AOI211_X1 g503(.A(KEYINPUT74), .B(new_n570), .C1(new_n583), .C2(new_n584), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n850), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n580), .A2(new_n624), .A3(new_n587), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n926), .B2(new_n932), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n925), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n925), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n867), .A2(new_n868), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n941), .ZN(G295));
  OAI21_X1  g517(.A(new_n940), .B1(G868), .B2(new_n941), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n551), .A2(new_n556), .B1(new_n867), .B2(new_n868), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n853), .A2(new_n854), .A3(new_n555), .A4(new_n858), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n945), .A2(G301), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(G286), .ZN(new_n949));
  OAI21_X1  g524(.A(G171), .B1(new_n859), .B2(new_n860), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(G301), .A3(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n934), .A3(new_n935), .ZN(new_n954));
  OAI21_X1  g529(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n931), .A3(new_n930), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n919), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n920), .A3(new_n958), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(KEYINPUT112), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT41), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT41), .B1(new_n930), .B2(new_n931), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n966), .A2(new_n957), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n953), .A2(new_n932), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n919), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n962), .ZN(new_n972));
  OR3_X1    g547(.A1(new_n972), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n944), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(KEYINPUT111), .A3(new_n963), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n977), .A3(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n974), .A2(new_n979), .ZN(G397));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n876), .B2(G1384), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT113), .B(G40), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n469), .A2(new_n478), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  INV_X1    g563(.A(new_n985), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n778), .B(new_n781), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(new_n764), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n764), .B(G1996), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n994), .A2(new_n990), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n829), .A2(new_n831), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n779), .A2(new_n781), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n989), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n829), .A2(new_n831), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1002), .A2(new_n985), .B1(KEYINPUT48), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1003), .A2(KEYINPUT48), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n999), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n993), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT127), .Z(new_n1008));
  NAND2_X1  g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n597), .A2(new_n598), .A3(new_n1011), .A4(new_n602), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n876), .A2(G1384), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n469), .A2(new_n478), .A3(new_n983), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n499), .A2(new_n496), .ZN(new_n1021));
  INV_X1    g596(.A(new_n875), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n874), .B1(new_n490), .B2(new_n493), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT115), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1013), .A2(new_n1014), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n591), .B(G1976), .C1(new_n594), .C2(new_n595), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1028), .B(new_n1030), .C1(new_n1019), .C2(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1015), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1025), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1033), .A2(new_n1034), .B1(G1976), .B2(new_n808), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1027), .B(new_n1031), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G166), .B2(new_n1016), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n984), .B1(new_n1017), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G164), .A2(G1384), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1045));
  INV_X1    g620(.A(new_n494), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1021), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1020), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1042), .A2(new_n1050), .A3(new_n732), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1024), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1018), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1971), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI221_X4 g631(.A(new_n1016), .B1(new_n1039), .B2(new_n1040), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(new_n876), .B2(G1384), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n732), .A4(new_n1018), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(KEYINPUT117), .A3(new_n1061), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G8), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(KEYINPUT118), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1042), .A2(new_n1050), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n707), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n982), .A2(new_n1018), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1048), .B2(new_n981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1044), .A2(KEYINPUT119), .A3(KEYINPUT45), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2078), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1054), .B2(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1072), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1069), .A2(new_n1070), .A3(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1075), .A2(new_n1076), .A3(new_n982), .A4(new_n1018), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n713), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1042), .A2(new_n1050), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT51), .B(G8), .C1(new_n1088), .C2(G286), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1016), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G168), .A2(new_n1016), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1091), .B(KEYINPUT51), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(G168), .B2(new_n1016), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1088), .A2(G8), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1097), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT124), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1090), .A2(new_n1094), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1102), .A2(KEYINPUT62), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT62), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1083), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1054), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1059), .A2(new_n1060), .A3(new_n1018), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n571), .B(new_n1114), .C1(new_n582), .C2(new_n581), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n585), .B2(new_n1114), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1348), .B1(new_n1042), .B2(new_n1050), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1025), .A2(G2067), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n624), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(KEYINPUT120), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT57), .B(new_n570), .C1(new_n573), .C2(new_n576), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(KEYINPUT57), .B2(new_n579), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT121), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1107), .A2(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1121), .A2(new_n1122), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1117), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n624), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n850), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1132), .B(new_n1136), .C1(KEYINPUT60), .C2(new_n1134), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1125), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1130), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1025), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1052), .A2(new_n986), .A3(new_n1018), .A4(new_n1053), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n557), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1144), .B2(new_n557), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT59), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1146), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1129), .B1(new_n1137), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1078), .A2(G40), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n982), .A2(new_n1052), .A3(G160), .A4(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1072), .A2(new_n1157), .A3(G301), .A4(new_n1080), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1069), .A2(new_n1070), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1072), .A2(new_n1080), .A3(new_n1157), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1072), .A2(new_n1079), .A3(G301), .A4(new_n1080), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(KEYINPUT54), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1163), .A2(KEYINPUT125), .A3(KEYINPUT54), .A4(new_n1164), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1155), .A2(new_n1160), .A3(new_n1161), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1064), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1172), .A2(new_n1062), .A3(new_n1016), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1173), .B2(new_n1066), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1099), .A2(G286), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1174), .A2(new_n1058), .A3(new_n1068), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1067), .B1(new_n1179), .B2(new_n1016), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1058), .A2(KEYINPUT63), .A3(new_n1175), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1057), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1037), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1027), .A2(new_n1029), .A3(new_n808), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1184), .A2(new_n1012), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT116), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1012), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT116), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1189), .B(new_n1190), .C1(new_n1182), .C2(new_n1037), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1178), .A2(new_n1181), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1106), .A2(new_n1170), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G290), .B(G1986), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n985), .B1(new_n1002), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1194), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1008), .B1(new_n1197), .B2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  OR4_X1    g775(.A1(new_n1201), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n905), .B2(new_n913), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n1203), .A2(new_n978), .A3(new_n976), .ZN(G308));
  NAND3_X1  g778(.A1(new_n1203), .A2(new_n978), .A3(new_n976), .ZN(G225));
endmodule


