//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n208), .A2(new_n210), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n221), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT86), .B(G50gat), .ZN(new_n223));
  INV_X1    g022(.A(G43gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n224), .A2(G50gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(new_n225), .B2(KEYINPUT87), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT15), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n220), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231));
  NAND2_X1  g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n231), .A2(new_n232), .B1(new_n233), .B2(KEYINPUT8), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT98), .B(G85gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(new_n235), .C1(G92gat), .C2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G99gat), .B(G106gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n230), .A2(new_n241), .B1(KEYINPUT41), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n205), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT99), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n244), .A3(new_n205), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n245), .B2(KEYINPUT99), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n203), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n245), .A2(KEYINPUT99), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(new_n246), .A3(new_n248), .A4(new_n202), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n243), .A2(KEYINPUT41), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT97), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n250), .B2(new_n252), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G183gat), .B(G211gat), .Z(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT96), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G71gat), .B(G78gat), .Z(new_n262));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT9), .ZN(new_n264));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G57gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G64gat), .ZN(new_n268));
  INV_X1    g067(.A(G64gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G57gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n264), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G71gat), .A2(G78gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT92), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n267), .B2(G64gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n269), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n268), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT94), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT94), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n282), .A4(new_n268), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n272), .B2(new_n264), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n276), .A2(KEYINPUT95), .A3(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT21), .ZN(new_n291));
  INV_X1    g090(.A(G231gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(G231gat), .B(G233gat), .C1(new_n290), .C2(KEYINPUT21), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n294), .B2(new_n295), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n261), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n297), .A3(new_n260), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT16), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n303), .A2(KEYINPUT88), .A3(G1gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT88), .B1(new_n303), .B2(G1gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G1gat), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT89), .B1(new_n305), .B2(G1gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G8gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n308), .B(new_n310), .Z(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n290), .B2(KEYINPUT21), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n300), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n300), .B2(new_n302), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n258), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n312), .ZN(new_n319));
  INV_X1    g118(.A(new_n258), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n257), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n288), .A2(new_n289), .A3(new_n239), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n239), .A2(new_n286), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n239), .A2(new_n327), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n290), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT100), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT100), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n324), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n325), .A2(new_n326), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n324), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G120gat), .B(G148gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G176gat), .B(G204gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n331), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n324), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n345), .B2(new_n338), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT101), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT101), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT90), .B1(new_n230), .B2(new_n240), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT90), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT17), .B1(new_n311), .B2(new_n354), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n353), .A2(new_n311), .B1(new_n355), .B2(new_n230), .ZN(new_n356));
  NAND2_X1  g155(.A1(G229gat), .A2(G233gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n230), .B(new_n311), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n357), .B(KEYINPUT13), .Z(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT18), .B1(new_n356), .B2(new_n357), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G141gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT11), .ZN(new_n366));
  INV_X1    g165(.A(G169gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G197gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT12), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n362), .A2(new_n363), .A3(new_n371), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT34), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n377), .A2(KEYINPUT65), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G183gat), .ZN(new_n380));
  INV_X1    g179(.A(G190gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT65), .B1(new_n377), .B2(new_n378), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n379), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT23), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(G169gat), .B2(G176gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n390), .B2(new_n387), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT25), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n378), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n382), .A3(new_n383), .ZN(new_n394));
  NAND2_X1  g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT23), .ZN(new_n396));
  OR2_X1    g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n398), .A2(new_n388), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT64), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n398), .B2(new_n388), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n394), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT28), .B1(new_n404), .B2(new_n381), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n380), .A2(KEYINPUT27), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT27), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G183gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT66), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n406), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n381), .A2(KEYINPUT28), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n405), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT26), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n397), .B2(KEYINPUT67), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n387), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n377), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n392), .B(new_n403), .C1(new_n415), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G113gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426));
  INV_X1    g225(.A(G120gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(G113gat), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(G113gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G134gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G127gat), .ZN(new_n432));
  INV_X1    g231(.A(G127gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G134gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n424), .A2(G120gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n434), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n430), .A2(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n391), .A2(KEYINPUT64), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n398), .A2(new_n388), .A3(new_n399), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n382), .B(new_n383), .C1(new_n393), .C2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n388), .B(new_n398), .C1(new_n446), .C2(new_n385), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n444), .A2(new_n394), .B1(new_n447), .B2(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n436), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n438), .A2(new_n439), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n377), .B(new_n421), .C1(new_n452), .C2(new_n405), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G227gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n293), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n376), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g258(.A(KEYINPUT34), .B(new_n457), .C1(new_n441), .C2(new_n454), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n457), .A3(new_n454), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT32), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G15gat), .B(G43gat), .Z(new_n466));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n462), .B(KEYINPUT32), .C1(new_n464), .C2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n461), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n459), .ZN(new_n473));
  INV_X1    g272(.A(new_n460), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n469), .A2(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT36), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n471), .ZN(new_n477));
  INV_X1    g276(.A(new_n461), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n469), .A3(new_n471), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G141gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(G148gat), .ZN(new_n487));
  INV_X1    g286(.A(G148gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(G141gat), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT71), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(G141gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(G148gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT2), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G155gat), .ZN(new_n498));
  INV_X1    g297(.A(G162gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n495), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n486), .A2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G141gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n505), .A3(G148gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n491), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n495), .B1(new_n500), .B2(KEYINPUT2), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n497), .A2(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT3), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G211gat), .B(G218gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G197gat), .B(G204gat), .ZN(new_n515));
  INV_X1    g314(.A(G211gat), .ZN(new_n516));
  INV_X1    g315(.A(G218gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n514), .B(new_n515), .C1(KEYINPUT22), .C2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G211gat), .B(G218gat), .Z(new_n520));
  INV_X1    g319(.A(G204gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G197gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n369), .A2(G204gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT22), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n519), .A2(new_n525), .A3(KEYINPUT69), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n494), .A2(new_n496), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n493), .B1(new_n491), .B2(new_n492), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n502), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n507), .A2(new_n508), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT29), .B1(new_n519), .B2(new_n525), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(KEYINPUT79), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n510), .B1(new_n538), .B2(KEYINPUT79), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G228gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n293), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n532), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n530), .B1(new_n511), .B2(new_n512), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n519), .B1(new_n525), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT78), .B1(new_n520), .B2(new_n524), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n512), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n509), .B1(new_n549), .B2(new_n510), .ZN(new_n550));
  OAI22_X1  g349(.A1(new_n545), .A2(new_n550), .B1(new_n542), .B2(new_n293), .ZN(new_n551));
  INV_X1    g350(.A(G22gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n544), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n544), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n485), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G22gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n544), .A2(new_n551), .A3(new_n552), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n484), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT31), .B(G50gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G226gat), .A2(G233gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n567), .B1(new_n423), .B2(new_n512), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n448), .B2(new_n453), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n568), .A2(new_n569), .A3(new_n531), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n531), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n574));
  OAI211_X1 g373(.A(KEYINPUT70), .B(new_n531), .C1(new_n568), .C2(new_n569), .ZN(new_n575));
  XNOR2_X1  g374(.A(G8gat), .B(G36gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G64gat), .B(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(new_n571), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n423), .A2(new_n512), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n566), .ZN(new_n583));
  INV_X1    g382(.A(new_n569), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n530), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n581), .A2(new_n575), .A3(new_n585), .A4(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT30), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n573), .B2(new_n575), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT4), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n440), .A2(new_n535), .A3(new_n590), .A4(new_n536), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n440), .A2(new_n535), .A3(new_n536), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n592), .A3(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n537), .A2(KEYINPUT3), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n511), .A3(new_n451), .ZN(new_n600));
  NAND2_X1  g399(.A1(G225gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT5), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n601), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n590), .A4(new_n440), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n608), .B1(KEYINPUT4), .B2(new_n594), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT74), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n509), .B2(new_n440), .ZN(new_n612));
  XNOR2_X1  g411(.A(G141gat), .B(G148gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n613), .A2(new_n493), .B1(KEYINPUT2), .B2(new_n495), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n501), .B1(new_n614), .B2(new_n490), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n501), .A2(new_n496), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n491), .B2(new_n506), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n451), .B(KEYINPUT74), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n612), .A2(new_n618), .B1(new_n509), .B2(new_n440), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT5), .B1(new_n619), .B2(new_n601), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n604), .B1(new_n610), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G1gat), .B(G29gat), .Z(new_n622));
  XNOR2_X1  g421(.A(G57gat), .B(G85gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n604), .B(new_n626), .C1(new_n610), .C2(new_n620), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n621), .A2(new_n627), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n589), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n483), .B1(new_n565), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n586), .A2(KEYINPUT30), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n586), .A2(KEYINPUT30), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n581), .A2(new_n575), .A3(new_n585), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n578), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n601), .B1(new_n598), .B2(new_n600), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n627), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n619), .B2(new_n601), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT80), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n440), .B1(new_n537), .B2(KEYINPUT3), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n596), .A2(new_n597), .B1(new_n511), .B2(new_n647), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n645), .A2(new_n646), .B1(new_n648), .B2(new_n601), .ZN(new_n649));
  INV_X1    g448(.A(new_n618), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT74), .B1(new_n537), .B2(new_n451), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n594), .B(new_n601), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n652), .A2(new_n646), .A3(KEYINPUT39), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n644), .B(KEYINPUT40), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  OAI221_X1 g453(.A(KEYINPUT5), .B1(new_n619), .B2(new_n601), .C1(new_n609), .C2(new_n605), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n626), .B1(new_n655), .B2(new_n604), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n644), .B1(new_n653), .B2(new_n649), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n641), .A2(KEYINPUT81), .A3(new_n654), .A4(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT81), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n646), .B1(new_n652), .B2(KEYINPUT39), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n653), .A2(new_n642), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n598), .A2(new_n600), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n643), .A3(new_n602), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n626), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n658), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n628), .A3(new_n654), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n668), .B2(new_n589), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n555), .A2(new_n559), .A3(new_n563), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n563), .B1(new_n555), .B2(new_n559), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n530), .B1(new_n583), .B2(new_n584), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT37), .B1(new_n674), .B2(new_n570), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n578), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT37), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n581), .A2(new_n678), .A3(new_n575), .A4(new_n585), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT82), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n573), .A2(KEYINPUT82), .A3(new_n678), .A4(new_n575), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n629), .A2(new_n631), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n633), .B(new_n586), .C1(new_n684), .C2(new_n656), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n579), .B1(new_n639), .B2(KEYINPUT37), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n676), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n673), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n636), .B1(new_n670), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT83), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT35), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n472), .A2(new_n475), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n562), .A2(new_n564), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(new_n635), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n640), .A2(KEYINPUT30), .A3(new_n586), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n697), .A2(new_n580), .B1(new_n632), .B2(new_n633), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n673), .A2(new_n698), .A3(KEYINPUT35), .A4(new_n694), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n691), .A2(new_n692), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n476), .A2(new_n482), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n698), .B2(new_n673), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n660), .A2(new_n669), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n688), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT38), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n683), .A2(new_n685), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n565), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT83), .B1(new_n710), .B2(new_n700), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n375), .B1(new_n702), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(KEYINPUT91), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT91), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n714), .B(new_n375), .C1(new_n702), .C2(new_n711), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n350), .B(new_n352), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n634), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT102), .B(G1gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1324gat));
  INV_X1    g518(.A(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n641), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n303), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n721), .A2(G8gat), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G8gat), .B1(new_n721), .B2(new_n724), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n722), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(G1325gat));
  OAI21_X1  g527(.A(G15gat), .B1(new_n716), .B2(new_n703), .ZN(new_n729));
  INV_X1    g528(.A(new_n694), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n730), .A2(G15gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n716), .B2(new_n731), .ZN(G1326gat));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n673), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  NAND2_X1  g534(.A1(new_n317), .A2(new_n321), .ZN(new_n736));
  INV_X1    g535(.A(new_n347), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n257), .ZN(new_n739));
  INV_X1    g538(.A(new_n375), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n692), .B1(new_n691), .B2(new_n701), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n710), .A2(KEYINPUT83), .A3(new_n700), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n714), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n712), .A2(KEYINPUT91), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n634), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n216), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n216), .A4(new_n747), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n691), .A2(KEYINPUT104), .A3(new_n701), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n710), .B2(new_n700), .ZN(new_n754));
  INV_X1    g553(.A(new_n257), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n702), .B2(new_n711), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n736), .A2(new_n375), .A3(new_n737), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n747), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n750), .B(new_n751), .C1(new_n216), .C2(new_n763), .ZN(G1328gat));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n217), .A3(new_n641), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n762), .A2(new_n641), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n767), .A2(new_n768), .B1(new_n217), .B2(new_n769), .ZN(G1329gat));
  AOI21_X1  g569(.A(G43gat), .B1(new_n746), .B2(new_n694), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n760), .A2(G43gat), .A3(new_n483), .A4(new_n761), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT106), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n777));
  INV_X1    g576(.A(new_n739), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n694), .B(new_n778), .C1(new_n713), .C2(new_n715), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n224), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(new_n781), .A3(new_n774), .A4(new_n772), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n776), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n777), .B1(new_n776), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1330gat));
  AOI21_X1  g584(.A(new_n223), .B1(new_n746), .B2(new_n565), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n565), .A2(new_n223), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n762), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1331gat));
  NAND3_X1  g589(.A1(new_n322), .A2(new_n375), .A3(new_n737), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT107), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n752), .A2(new_n754), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n634), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n267), .ZN(G1332gat));
  INV_X1    g595(.A(new_n794), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n641), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n799), .B2(new_n798), .ZN(G1333gat));
  NAND3_X1  g601(.A1(new_n797), .A2(G71gat), .A3(new_n483), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G71gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n794), .B2(new_n730), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n797), .A2(new_n565), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g611(.A1(new_n317), .A2(new_n321), .A3(new_n257), .A4(new_n375), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n691), .B2(new_n701), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT109), .B1(new_n814), .B2(KEYINPUT51), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n710), .A2(new_n700), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(new_n813), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(KEYINPUT51), .C1(new_n710), .C2(new_n700), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n737), .ZN(new_n823));
  INV_X1    g622(.A(new_n236), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n747), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n736), .A2(new_n740), .A3(new_n347), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n760), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n236), .B1(new_n827), .B2(new_n634), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1336gat));
  INV_X1    g628(.A(G92gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n702), .A2(new_n711), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n759), .B1(new_n831), .B2(new_n257), .ZN(new_n832));
  INV_X1    g631(.A(new_n757), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n641), .B(new_n826), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n641), .A4(new_n826), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n347), .A2(G92gat), .A3(new_n589), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT111), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT111), .B1(new_n822), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n691), .A2(new_n701), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(new_n845), .B2(new_n820), .ZN(new_n846));
  INV_X1    g645(.A(new_n821), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n840), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT110), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n840), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(G92gat), .B2(new_n834), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n838), .A2(new_n844), .B1(new_n853), .B2(new_n839), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n834), .A2(G92gat), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT52), .B1(new_n856), .B2(new_n852), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n857), .B(new_n858), .C1(new_n838), .C2(new_n844), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(G1337gat));
  INV_X1    g659(.A(G99gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n823), .A2(new_n861), .A3(new_n694), .ZN(new_n862));
  OAI21_X1  g661(.A(G99gat), .B1(new_n827), .B2(new_n703), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1338gat));
  INV_X1    g663(.A(G106gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n823), .A2(new_n865), .A3(new_n565), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n760), .A2(new_n565), .A3(new_n826), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT114), .B(G106gat), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n846), .A2(new_n847), .ZN(new_n874));
  NOR4_X1   g673(.A1(new_n874), .A2(G106gat), .A3(new_n673), .A4(new_n347), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT53), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n872), .B1(new_n868), .B2(new_n871), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(G1339gat));
  NOR2_X1   g677(.A1(new_n641), .A2(new_n634), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n736), .ZN(new_n881));
  INV_X1    g680(.A(new_n334), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n333), .B1(new_n328), .B2(new_n330), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n323), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT54), .B1(new_n331), .B2(new_n323), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(KEYINPUT116), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n341), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n345), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n335), .B2(new_n885), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n887), .A3(KEYINPUT55), .A4(new_n890), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n893), .A2(new_n887), .A3(new_n890), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n342), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n740), .A3(new_n901), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n356), .A2(new_n357), .B1(new_n360), .B2(new_n359), .ZN(new_n903));
  INV_X1    g702(.A(new_n370), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n374), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n347), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n257), .B1(new_n902), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n907), .A2(new_n255), .A3(new_n256), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n898), .A3(new_n901), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n881), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n348), .A2(new_n740), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n880), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n695), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n740), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n737), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(KEYINPUT118), .A3(new_n427), .ZN(new_n923));
  XNOR2_X1  g722(.A(KEYINPUT118), .B(G120gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(G1341gat));
  NAND2_X1  g724(.A1(new_n919), .A2(new_n736), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g726(.A1(new_n919), .A2(new_n257), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G134gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n919), .A2(new_n431), .A3(new_n257), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT119), .B1(new_n930), .B2(KEYINPUT56), .ZN(new_n932));
  OAI221_X1 g731(.A(new_n929), .B1(KEYINPUT56), .B2(new_n930), .C1(new_n931), .C2(new_n932), .ZN(G1343gat));
  NOR2_X1   g732(.A1(new_n673), .A2(new_n483), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n917), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(new_n486), .A3(new_n740), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT58), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n503), .A2(new_n505), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n880), .A2(new_n483), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n914), .A2(new_n916), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n940), .B2(new_n565), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n343), .B1(new_n373), .B2(new_n374), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n897), .B2(new_n894), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n900), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n908), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n912), .B1(new_n947), .B2(new_n257), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n915), .B1(new_n948), .B2(new_n881), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n565), .A2(KEYINPUT57), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n939), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n938), .B1(new_n952), .B2(new_n375), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(KEYINPUT121), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n673), .B1(new_n914), .B2(new_n916), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n956), .A2(KEYINPUT57), .B1(new_n949), .B2(new_n950), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n958), .A3(new_n939), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n740), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n936), .B1(new_n960), .B2(new_n938), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT58), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n954), .B1(new_n961), .B2(new_n962), .ZN(G1344gat));
  AND3_X1   g762(.A1(new_n957), .A2(new_n958), .A3(new_n939), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n958), .B1(new_n957), .B2(new_n939), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n964), .A2(new_n965), .A3(new_n347), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G148gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT57), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n956), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n565), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n352), .A2(new_n375), .A3(new_n350), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n881), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n970), .A2(new_n974), .A3(new_n347), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n488), .B1(new_n975), .B2(new_n939), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n966), .A2(new_n968), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NOR4_X1   g776(.A1(new_n347), .A2(new_n641), .A3(G148gat), .A4(new_n634), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n940), .A2(new_n934), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1345gat));
  AOI21_X1  g779(.A(G155gat), .B1(new_n935), .B2(new_n736), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n965), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n736), .A2(G155gat), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT122), .Z(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n982), .B2(new_n984), .ZN(G1346gat));
  NAND3_X1  g784(.A1(new_n935), .A2(new_n499), .A3(new_n257), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n964), .A2(new_n965), .A3(new_n755), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n499), .ZN(G1347gat));
  AOI21_X1  g787(.A(new_n747), .B1(new_n914), .B2(new_n916), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(new_n641), .A3(new_n918), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n740), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n737), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(G176gat), .ZN(G1349gat));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n990), .A2(new_n412), .A3(new_n736), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n990), .A2(new_n736), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n995), .B(new_n996), .C1(new_n997), .C2(new_n380), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g798(.A1(new_n990), .A2(new_n257), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G190gat), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT61), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1002), .B1(G190gat), .B2(new_n1000), .ZN(G1351gat));
  NAND2_X1  g802(.A1(new_n934), .A2(new_n641), .ZN(new_n1004));
  XOR2_X1   g803(.A(new_n1004), .B(KEYINPUT124), .Z(new_n1005));
  AND2_X1   g804(.A1(new_n989), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g805(.A(KEYINPUT125), .B(G197gat), .Z(new_n1007));
  NAND3_X1  g806(.A1(new_n1006), .A2(new_n740), .A3(new_n1007), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n483), .A2(new_n747), .A3(new_n589), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n970), .A2(new_n974), .A3(new_n1010), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1011), .A2(new_n740), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1008), .B1(new_n1012), .B2(new_n1007), .ZN(G1352gat));
  AOI21_X1  g812(.A(new_n521), .B1(new_n975), .B2(new_n1009), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n347), .A2(G204gat), .ZN(new_n1017));
  NAND4_X1  g816(.A1(new_n989), .A2(new_n1016), .A3(new_n1005), .A4(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT126), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n1015), .A2(KEYINPUT127), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1023), .B1(new_n1024), .B2(new_n1014), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1022), .A2(new_n1025), .ZN(G1353gat));
  NAND3_X1  g825(.A1(new_n1006), .A2(new_n516), .A3(new_n736), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n736), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n1028), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1029));
  AOI21_X1  g828(.A(KEYINPUT63), .B1(new_n1028), .B2(G211gat), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G1354gat));
  NAND3_X1  g830(.A1(new_n1006), .A2(new_n517), .A3(new_n257), .ZN(new_n1032));
  AND2_X1   g831(.A1(new_n1011), .A2(new_n257), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1032), .B1(new_n1033), .B2(new_n517), .ZN(G1355gat));
endmodule


