

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n599), .A2(n598), .ZN(n1009) );
  XNOR2_X1 U555 ( .A(n597), .B(KEYINPUT72), .ZN(n599) );
  XNOR2_X2 U556 ( .A(n798), .B(KEYINPUT103), .ZN(n799) );
  AND2_X2 U557 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U558 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U559 ( .A1(n702), .A2(n819), .ZN(n758) );
  XNOR2_X1 U560 ( .A(KEYINPUT91), .B(n818), .ZN(n702) );
  BUF_X1 U561 ( .A(n624), .Z(n625) );
  NOR2_X2 U562 ( .A1(G2104), .A2(n522), .ZN(n911) );
  XNOR2_X1 U563 ( .A(KEYINPUT94), .B(n729), .ZN(n733) );
  INV_X1 U564 ( .A(KEYINPUT97), .ZN(n722) );
  AND2_X1 U565 ( .A1(n717), .A2(n710), .ZN(n711) );
  INV_X1 U566 ( .A(n758), .ZN(n724) );
  BUF_X1 U567 ( .A(n724), .Z(n738) );
  XNOR2_X1 U568 ( .A(n767), .B(KEYINPUT100), .ZN(n768) );
  INV_X1 U569 ( .A(n778), .ZN(n779) );
  NAND2_X1 U570 ( .A1(n780), .A2(n779), .ZN(n781) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n904), .A2(n527), .ZN(n530) );
  NAND2_X1 U573 ( .A1(n831), .A2(n840), .ZN(n832) );
  OR2_X1 U574 ( .A1(n833), .A2(n832), .ZN(n847) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X2 U576 ( .A(n519), .B(n518), .ZN(n904) );
  NAND2_X1 U577 ( .A1(G138), .A2(n904), .ZN(n521) );
  INV_X1 U578 ( .A(G2105), .ZN(n522) );
  AND2_X1 U579 ( .A1(n522), .A2(G2104), .ZN(n624) );
  NAND2_X1 U580 ( .A1(G102), .A2(n624), .ZN(n520) );
  NAND2_X1 U581 ( .A1(n521), .A2(n520), .ZN(n526) );
  NAND2_X1 U582 ( .A1(G126), .A2(n911), .ZN(n524) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n908) );
  NAND2_X1 U584 ( .A1(G114), .A2(n908), .ZN(n523) );
  NAND2_X1 U585 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U586 ( .A1(n526), .A2(n525), .ZN(G164) );
  AND2_X1 U587 ( .A1(G137), .A2(KEYINPUT65), .ZN(n527) );
  INV_X1 U588 ( .A(KEYINPUT65), .ZN(n528) );
  NAND2_X1 U589 ( .A1(G113), .A2(n908), .ZN(n531) );
  OR2_X1 U590 ( .A1(n528), .A2(n531), .ZN(n529) );
  AND2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n904), .A2(G137), .ZN(n533) );
  AND2_X1 U593 ( .A1(n528), .A2(n531), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n701) );
  NAND2_X1 U596 ( .A1(G101), .A2(n624), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT23), .ZN(n538) );
  INV_X1 U598 ( .A(KEYINPUT64), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n538), .B(n537), .ZN(n699) );
  NAND2_X1 U600 ( .A1(G125), .A2(n911), .ZN(n697) );
  AND2_X1 U601 ( .A1(n699), .A2(n697), .ZN(n539) );
  AND2_X1 U602 ( .A1(n701), .A2(n539), .ZN(G160) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n667) );
  INV_X1 U604 ( .A(G651), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n667), .A2(n542), .ZN(n650) );
  NAND2_X1 U606 ( .A1(G78), .A2(n650), .ZN(n541) );
  NOR2_X2 U607 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U608 ( .A1(G91), .A2(n652), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n547) );
  NOR2_X1 U610 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT1), .B(n543), .Z(n592) );
  BUF_X1 U612 ( .A(n592), .Z(n663) );
  NAND2_X1 U613 ( .A1(G65), .A2(n663), .ZN(n545) );
  NOR2_X2 U614 ( .A1(n667), .A2(G651), .ZN(n660) );
  NAND2_X1 U615 ( .A1(G53), .A2(n660), .ZN(n544) );
  NAND2_X1 U616 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U617 ( .A1(n547), .A2(n546), .ZN(G299) );
  XOR2_X1 U618 ( .A(G2443), .B(G2446), .Z(n549) );
  XNOR2_X1 U619 ( .A(G2427), .B(G2451), .ZN(n548) );
  XNOR2_X1 U620 ( .A(n549), .B(n548), .ZN(n555) );
  XOR2_X1 U621 ( .A(G2430), .B(G2454), .Z(n551) );
  XNOR2_X1 U622 ( .A(G1341), .B(G1348), .ZN(n550) );
  XNOR2_X1 U623 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U624 ( .A(G2435), .B(G2438), .Z(n552) );
  XNOR2_X1 U625 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U626 ( .A(n555), .B(n554), .Z(n556) );
  AND2_X1 U627 ( .A1(G14), .A2(n556), .ZN(G401) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(n650), .A2(G75), .ZN(n559) );
  NAND2_X1 U633 ( .A1(G88), .A2(n652), .ZN(n557) );
  XOR2_X1 U634 ( .A(KEYINPUT83), .B(n557), .Z(n558) );
  NAND2_X1 U635 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U636 ( .A1(G62), .A2(n663), .ZN(n561) );
  NAND2_X1 U637 ( .A1(G50), .A2(n660), .ZN(n560) );
  NAND2_X1 U638 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U639 ( .A1(n563), .A2(n562), .ZN(G166) );
  XNOR2_X1 U640 ( .A(KEYINPUT69), .B(KEYINPUT9), .ZN(n567) );
  NAND2_X1 U641 ( .A1(G77), .A2(n650), .ZN(n565) );
  NAND2_X1 U642 ( .A1(G90), .A2(n652), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U644 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n663), .A2(G64), .ZN(n568) );
  XNOR2_X1 U646 ( .A(n568), .B(KEYINPUT68), .ZN(n570) );
  NAND2_X1 U647 ( .A1(G52), .A2(n660), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U649 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U650 ( .A1(n652), .A2(G89), .ZN(n573) );
  XNOR2_X1 U651 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U652 ( .A1(G76), .A2(n650), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U654 ( .A(KEYINPUT5), .B(n576), .ZN(n583) );
  XNOR2_X1 U655 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G63), .A2(n663), .ZN(n578) );
  NAND2_X1 U657 ( .A1(G51), .A2(n660), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U659 ( .A(n579), .B(KEYINPUT6), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n581), .B(n580), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U662 ( .A(KEYINPUT7), .B(n584), .ZN(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT10), .ZN(n586) );
  XNOR2_X1 U666 ( .A(KEYINPUT70), .B(n586), .ZN(G223) );
  INV_X1 U667 ( .A(G223), .ZN(n849) );
  NAND2_X1 U668 ( .A1(n849), .A2(G567), .ZN(n587) );
  XOR2_X1 U669 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U670 ( .A1(n652), .A2(G81), .ZN(n588) );
  XNOR2_X1 U671 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n650), .A2(G68), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U674 ( .A(KEYINPUT13), .B(n591), .Z(n596) );
  NAND2_X1 U675 ( .A1(G56), .A2(n592), .ZN(n593) );
  XNOR2_X1 U676 ( .A(n593), .B(KEYINPUT71), .ZN(n594) );
  XNOR2_X1 U677 ( .A(n594), .B(KEYINPUT14), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U679 ( .A1(G43), .A2(n660), .ZN(n598) );
  INV_X1 U680 ( .A(G860), .ZN(n614) );
  OR2_X1 U681 ( .A1(n1009), .A2(n614), .ZN(G153) );
  INV_X1 U682 ( .A(G171), .ZN(G301) );
  NAND2_X1 U683 ( .A1(G66), .A2(n663), .ZN(n606) );
  NAND2_X1 U684 ( .A1(G79), .A2(n650), .ZN(n601) );
  NAND2_X1 U685 ( .A1(G92), .A2(n652), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U687 ( .A1(G54), .A2(n660), .ZN(n602) );
  XNOR2_X1 U688 ( .A(KEYINPUT73), .B(n602), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(KEYINPUT15), .ZN(n608) );
  XOR2_X1 U692 ( .A(KEYINPUT74), .B(n608), .Z(n709) );
  BUF_X1 U693 ( .A(n709), .Z(n1022) );
  NOR2_X1 U694 ( .A1(n1022), .A2(G868), .ZN(n610) );
  INV_X1 U695 ( .A(G868), .ZN(n670) );
  NOR2_X1 U696 ( .A1(n670), .A2(G301), .ZN(n609) );
  NOR2_X1 U697 ( .A1(n610), .A2(n609), .ZN(G284) );
  NOR2_X1 U698 ( .A1(G286), .A2(n670), .ZN(n612) );
  NOR2_X1 U699 ( .A1(G868), .A2(G299), .ZN(n611) );
  NOR2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U701 ( .A(KEYINPUT77), .B(n613), .Z(G297) );
  NAND2_X1 U702 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U703 ( .A(n615), .B(KEYINPUT78), .ZN(n616) );
  INV_X1 U704 ( .A(n1022), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n616), .A2(n632), .ZN(n617) );
  XNOR2_X1 U706 ( .A(KEYINPUT16), .B(n617), .ZN(G148) );
  NOR2_X1 U707 ( .A1(G868), .A2(n1009), .ZN(n620) );
  NAND2_X1 U708 ( .A1(n632), .A2(G868), .ZN(n618) );
  NOR2_X1 U709 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U710 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U711 ( .A1(n911), .A2(G123), .ZN(n621) );
  XNOR2_X1 U712 ( .A(n621), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U713 ( .A1(G111), .A2(n908), .ZN(n622) );
  NAND2_X1 U714 ( .A1(n623), .A2(n622), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G135), .A2(n904), .ZN(n627) );
  NAND2_X1 U716 ( .A1(G99), .A2(n625), .ZN(n626) );
  NAND2_X1 U717 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n935) );
  XNOR2_X1 U719 ( .A(n935), .B(G2096), .ZN(n631) );
  INV_X1 U720 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U721 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U722 ( .A1(n632), .A2(G559), .ZN(n633) );
  XNOR2_X1 U723 ( .A(n633), .B(n1009), .ZN(n679) );
  NOR2_X1 U724 ( .A1(n679), .A2(G860), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G67), .A2(n663), .ZN(n635) );
  NAND2_X1 U726 ( .A1(G55), .A2(n660), .ZN(n634) );
  NAND2_X1 U727 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U728 ( .A1(G80), .A2(n650), .ZN(n636) );
  XNOR2_X1 U729 ( .A(KEYINPUT79), .B(n636), .ZN(n637) );
  NOR2_X1 U730 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n652), .A2(G93), .ZN(n639) );
  NAND2_X1 U732 ( .A1(n640), .A2(n639), .ZN(n672) );
  XOR2_X1 U733 ( .A(n641), .B(n672), .Z(G145) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n643) );
  NAND2_X1 U735 ( .A1(G73), .A2(n650), .ZN(n642) );
  XNOR2_X1 U736 ( .A(n643), .B(n642), .ZN(n647) );
  NAND2_X1 U737 ( .A1(G86), .A2(n652), .ZN(n645) );
  NAND2_X1 U738 ( .A1(G61), .A2(n663), .ZN(n644) );
  NAND2_X1 U739 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U740 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n660), .A2(G48), .ZN(n648) );
  NAND2_X1 U742 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U743 ( .A1(n650), .A2(G72), .ZN(n651) );
  XNOR2_X1 U744 ( .A(n651), .B(KEYINPUT66), .ZN(n654) );
  NAND2_X1 U745 ( .A1(G85), .A2(n652), .ZN(n653) );
  NAND2_X1 U746 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U747 ( .A(KEYINPUT67), .B(n655), .ZN(n659) );
  NAND2_X1 U748 ( .A1(G60), .A2(n663), .ZN(n657) );
  NAND2_X1 U749 ( .A1(G47), .A2(n660), .ZN(n656) );
  AND2_X1 U750 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U751 ( .A1(n659), .A2(n658), .ZN(G290) );
  NAND2_X1 U752 ( .A1(n660), .A2(G49), .ZN(n661) );
  XOR2_X1 U753 ( .A(KEYINPUT80), .B(n661), .Z(n662) );
  NOR2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U755 ( .A1(G651), .A2(G74), .ZN(n664) );
  NAND2_X1 U756 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U757 ( .A(n666), .B(KEYINPUT81), .ZN(n669) );
  NAND2_X1 U758 ( .A1(G87), .A2(n667), .ZN(n668) );
  NAND2_X1 U759 ( .A1(n669), .A2(n668), .ZN(G288) );
  AND2_X1 U760 ( .A1(n670), .A2(n672), .ZN(n671) );
  XNOR2_X1 U761 ( .A(n671), .B(KEYINPUT85), .ZN(n682) );
  XNOR2_X1 U762 ( .A(KEYINPUT19), .B(G299), .ZN(n673) );
  XNOR2_X1 U763 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U764 ( .A(KEYINPUT84), .B(n674), .ZN(n676) );
  XNOR2_X1 U765 ( .A(G305), .B(G166), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U767 ( .A(n677), .B(G290), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(G288), .ZN(n919) );
  XNOR2_X1 U769 ( .A(n919), .B(n679), .ZN(n680) );
  NAND2_X1 U770 ( .A1(G868), .A2(n680), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(G295) );
  NAND2_X1 U772 ( .A1(G2078), .A2(G2084), .ZN(n683) );
  XOR2_X1 U773 ( .A(KEYINPUT20), .B(n683), .Z(n684) );
  NAND2_X1 U774 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U775 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U777 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U778 ( .A1(G120), .A2(G69), .ZN(n687) );
  NOR2_X1 U779 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U780 ( .A1(G108), .A2(n688), .ZN(n856) );
  NAND2_X1 U781 ( .A1(n856), .A2(G567), .ZN(n694) );
  NOR2_X1 U782 ( .A1(G220), .A2(G219), .ZN(n689) );
  XOR2_X1 U783 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U784 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U785 ( .A1(G96), .A2(n691), .ZN(n855) );
  NAND2_X1 U786 ( .A1(G2106), .A2(n855), .ZN(n692) );
  XNOR2_X1 U787 ( .A(KEYINPUT86), .B(n692), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n932) );
  NAND2_X1 U789 ( .A1(G661), .A2(G483), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT87), .B(n695), .Z(n696) );
  NOR2_X1 U791 ( .A1(n932), .A2(n696), .ZN(n854) );
  NAND2_X1 U792 ( .A1(n854), .A2(G36), .ZN(G176) );
  INV_X1 U793 ( .A(G166), .ZN(G303) );
  AND2_X1 U794 ( .A1(n697), .A2(G40), .ZN(n698) );
  AND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n818) );
  NOR2_X1 U797 ( .A1(G164), .A2(G1384), .ZN(n819) );
  NAND2_X1 U798 ( .A1(G8), .A2(n758), .ZN(n778) );
  NOR2_X1 U799 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U800 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  NOR2_X1 U801 ( .A1(n778), .A2(n704), .ZN(n800) );
  NOR2_X1 U802 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n758), .ZN(n744) );
  NAND2_X1 U804 ( .A1(n744), .A2(G8), .ZN(n755) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n778), .ZN(n753) );
  INV_X1 U806 ( .A(KEYINPUT26), .ZN(n706) );
  NAND2_X1 U807 ( .A1(G1996), .A2(n724), .ZN(n705) );
  XNOR2_X1 U808 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X2 U809 ( .A1(n707), .A2(n1009), .ZN(n717) );
  NAND2_X1 U810 ( .A1(G1341), .A2(n758), .ZN(n718) );
  INV_X1 U811 ( .A(n718), .ZN(n708) );
  NOR2_X1 U812 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U813 ( .A(n711), .B(KEYINPUT95), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n758), .A2(G1348), .ZN(n712) );
  XNOR2_X1 U815 ( .A(n712), .B(KEYINPUT96), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n738), .A2(G2067), .ZN(n713) );
  NAND2_X1 U817 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n717), .A2(n718), .ZN(n719) );
  NAND2_X1 U820 ( .A1(n1022), .A2(n719), .ZN(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U822 ( .A(n723), .B(n722), .ZN(n732) );
  AND2_X1 U823 ( .A1(n724), .A2(G2072), .ZN(n726) );
  XNOR2_X1 U824 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n725) );
  XNOR2_X1 U825 ( .A(n726), .B(n725), .ZN(n728) );
  XOR2_X1 U826 ( .A(KEYINPUT93), .B(G1956), .Z(n961) );
  NAND2_X1 U827 ( .A1(n758), .A2(n961), .ZN(n727) );
  NAND2_X1 U828 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U829 ( .A1(n733), .A2(G299), .ZN(n730) );
  XOR2_X1 U830 ( .A(KEYINPUT98), .B(n730), .Z(n731) );
  NAND2_X1 U831 ( .A1(n732), .A2(n731), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n733), .A2(G299), .ZN(n734) );
  XNOR2_X1 U833 ( .A(n734), .B(KEYINPUT28), .ZN(n735) );
  NAND2_X1 U834 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U835 ( .A(n737), .B(KEYINPUT29), .ZN(n742) );
  XOR2_X1 U836 ( .A(G2078), .B(KEYINPUT25), .Z(n994) );
  NOR2_X1 U837 ( .A1(n994), .A2(n758), .ZN(n740) );
  NOR2_X1 U838 ( .A1(n738), .A2(G1961), .ZN(n739) );
  NOR2_X1 U839 ( .A1(n740), .A2(n739), .ZN(n743) );
  NOR2_X1 U840 ( .A1(G301), .A2(n743), .ZN(n741) );
  NOR2_X1 U841 ( .A1(n742), .A2(n741), .ZN(n752) );
  AND2_X1 U842 ( .A1(G301), .A2(n743), .ZN(n749) );
  NOR2_X1 U843 ( .A1(n753), .A2(n744), .ZN(n745) );
  NAND2_X1 U844 ( .A1(G8), .A2(n745), .ZN(n746) );
  XNOR2_X1 U845 ( .A(KEYINPUT30), .B(n746), .ZN(n747) );
  NOR2_X1 U846 ( .A1(G168), .A2(n747), .ZN(n748) );
  NOR2_X1 U847 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U848 ( .A(n750), .B(KEYINPUT31), .ZN(n751) );
  NOR2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n753), .A2(n757), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n771) );
  INV_X1 U852 ( .A(G286), .ZN(n756) );
  OR2_X1 U853 ( .A1(n757), .A2(n756), .ZN(n766) );
  INV_X1 U854 ( .A(G8), .ZN(n764) );
  NOR2_X1 U855 ( .A1(G1971), .A2(n778), .ZN(n760) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U858 ( .A(KEYINPUT99), .B(n761), .Z(n762) );
  NAND2_X1 U859 ( .A1(n762), .A2(G303), .ZN(n763) );
  OR2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U861 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n767) );
  XNOR2_X1 U862 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n783) );
  INV_X1 U864 ( .A(G1971), .ZN(n975) );
  NAND2_X1 U865 ( .A1(G166), .A2(n975), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n783), .A2(n772), .ZN(n773) );
  NOR2_X1 U867 ( .A1(n1015), .A2(n773), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n1025) );
  INV_X1 U869 ( .A(KEYINPUT33), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n779), .A2(n1015), .ZN(n774) );
  NOR2_X1 U871 ( .A1(n786), .A2(n774), .ZN(n775) );
  XOR2_X1 U872 ( .A(n775), .B(KEYINPUT102), .Z(n785) );
  AND2_X1 U873 ( .A1(n1025), .A2(n785), .ZN(n777) );
  XNOR2_X1 U874 ( .A(G1981), .B(G305), .ZN(n1011) );
  INV_X1 U875 ( .A(n1011), .ZN(n776) );
  AND2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n780) );
  OR2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n797) );
  INV_X1 U878 ( .A(n783), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G8), .A2(G166), .ZN(n784) );
  NOR2_X1 U880 ( .A1(G2090), .A2(n784), .ZN(n790) );
  INV_X1 U881 ( .A(n785), .ZN(n787) );
  OR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U883 ( .A1(n1011), .A2(n788), .ZN(n793) );
  INV_X1 U884 ( .A(n793), .ZN(n789) );
  OR2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n795) );
  AND2_X1 U887 ( .A1(n793), .A2(n779), .ZN(n794) );
  OR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n833) );
  XOR2_X1 U890 ( .A(G1986), .B(G290), .Z(n1016) );
  NAND2_X1 U891 ( .A1(G131), .A2(n904), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G119), .A2(n911), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G95), .A2(n625), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G107), .A2(n908), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n897) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n897), .ZN(n816) );
  NAND2_X1 U899 ( .A1(G141), .A2(n904), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G129), .A2(n911), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G105), .A2(n625), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT38), .ZN(n810) );
  XNOR2_X1 U904 ( .A(n810), .B(KEYINPUT89), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n908), .A2(G117), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n886) );
  NAND2_X1 U908 ( .A1(G1996), .A2(n886), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U910 ( .A(KEYINPUT90), .B(n817), .Z(n834) );
  NAND2_X1 U911 ( .A1(n1016), .A2(n834), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n844) );
  NAND2_X1 U913 ( .A1(n820), .A2(n844), .ZN(n831) );
  XNOR2_X1 U914 ( .A(KEYINPUT37), .B(G2067), .ZN(n842) );
  NAND2_X1 U915 ( .A1(G140), .A2(n904), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G104), .A2(n625), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U918 ( .A(KEYINPUT34), .B(n823), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G128), .A2(n911), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G116), .A2(n908), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT88), .B(n826), .Z(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT35), .B(n827), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT36), .B(n830), .ZN(n901) );
  NOR2_X1 U926 ( .A1(n842), .A2(n901), .ZN(n934) );
  NAND2_X1 U927 ( .A1(n844), .A2(n934), .ZN(n840) );
  INV_X1 U928 ( .A(n834), .ZN(n940) );
  NOR2_X1 U929 ( .A1(G1991), .A2(n897), .ZN(n936) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n936), .A2(n835), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n940), .A2(n836), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n886), .A2(G1996), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n837), .B(KEYINPUT104), .ZN(n949) );
  NOR2_X1 U935 ( .A1(n838), .A2(n949), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT39), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n842), .A2(n901), .ZN(n937) );
  NAND2_X1 U939 ( .A1(n843), .A2(n937), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U942 ( .A(n848), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n849), .ZN(G217) );
  NAND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n851) );
  INV_X1 U945 ( .A(G661), .ZN(n850) );
  NOR2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(G188) );
  XOR2_X1 U950 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G325) );
  XNOR2_X1 U952 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U954 ( .A(G120), .ZN(G236) );
  INV_X1 U955 ( .A(G96), .ZN(G221) );
  XOR2_X1 U956 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2072), .B(KEYINPUT108), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n859), .B(G2678), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2090), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT42), .B(G2100), .Z(n863) );
  XNOR2_X1 U963 ( .A(G2078), .B(G2084), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G227) );
  XOR2_X1 U966 ( .A(G1966), .B(G1956), .Z(n867) );
  XNOR2_X1 U967 ( .A(G1981), .B(G1971), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n877) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1991), .B(KEYINPUT111), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U972 ( .A(G1976), .B(G1961), .Z(n871) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1986), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U976 ( .A(KEYINPUT110), .B(G2474), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(n877), .B(n876), .Z(G229) );
  NAND2_X1 U979 ( .A1(n911), .A2(G124), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G112), .A2(n908), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G136), .A2(n904), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G100), .A2(n625), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U987 ( .A(G164), .B(G162), .Z(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n935), .B(n887), .ZN(n903) );
  XNOR2_X1 U990 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n899) );
  NAND2_X1 U991 ( .A1(n904), .A2(G139), .ZN(n888) );
  XNOR2_X1 U992 ( .A(KEYINPUT113), .B(n888), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G127), .A2(n911), .ZN(n890) );
  NAND2_X1 U994 ( .A1(G115), .A2(n908), .ZN(n889) );
  NAND2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n891), .B(KEYINPUT114), .ZN(n892) );
  XNOR2_X1 U997 ( .A(n892), .B(KEYINPUT47), .ZN(n894) );
  NAND2_X1 U998 ( .A1(n625), .A2(G103), .ZN(n893) );
  NAND2_X1 U999 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U1000 ( .A1(n896), .A2(n895), .ZN(n944) );
  XNOR2_X1 U1001 ( .A(n897), .B(n944), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1003 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n917) );
  NAND2_X1 U1005 ( .A1(G142), .A2(n904), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(G106), .A2(n625), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n907), .B(KEYINPUT45), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(G118), .A2(n908), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n911), .A2(G130), .ZN(n912) );
  XOR2_X1 U1012 ( .A(KEYINPUT112), .B(n912), .Z(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(G160), .B(n915), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1017 ( .A(KEYINPUT115), .B(n919), .Z(n921) );
  XNOR2_X1 U1018 ( .A(G171), .B(n1022), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n921), .B(n920), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n1009), .B(G286), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n924), .ZN(G397) );
  NOR2_X1 U1023 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT49), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT117), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G401), .A2(n932), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n929), .B(KEYINPUT116), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(n932), .ZN(G319) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1034 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n955) );
  XNOR2_X1 U1040 ( .A(G164), .B(G2078), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(n943), .B(KEYINPUT119), .ZN(n946) );
  XOR2_X1 U1042 ( .A(n944), .B(G2072), .Z(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT50), .B(n947), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1047 ( .A(KEYINPUT118), .B(n950), .Z(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT51), .B(n951), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT52), .B(n956), .ZN(n958) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(G29), .ZN(n1038) );
  XOR2_X1 U1055 ( .A(G1961), .B(G5), .Z(n974) );
  XOR2_X1 U1056 ( .A(G1348), .B(KEYINPUT59), .Z(n960) );
  XNOR2_X1 U1057 ( .A(G4), .B(n960), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G20), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1981), .B(G6), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G19), .B(G1341), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT60), .ZN(n969) );
  XOR2_X1 U1065 ( .A(KEYINPUT125), .B(n969), .Z(n971) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT126), .B(n972), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n982) );
  XOR2_X1 U1070 ( .A(G1986), .B(G24), .Z(n977) );
  XNOR2_X1 U1071 ( .A(n975), .B(G22), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G23), .B(G1976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1075 ( .A(KEYINPUT58), .B(n980), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n983), .Z(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT124), .B(G16), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n1036) );
  XNOR2_X1 U1080 ( .A(G1996), .B(G32), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G33), .B(G2072), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n993) );
  XOR2_X1 U1083 ( .A(G2067), .B(G26), .Z(n988) );
  NAND2_X1 U1084 ( .A1(n988), .A2(G28), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(G25), .B(G1991), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(KEYINPUT120), .B(n989), .ZN(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G27), .B(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1091 ( .A(KEYINPUT53), .B(n997), .Z(n1000) );
  XOR2_X1 U1092 ( .A(G34), .B(KEYINPUT54), .Z(n998) );
  XNOR2_X1 U1093 ( .A(G2084), .B(n998), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(G35), .B(G2090), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1097 ( .A(KEYINPUT55), .B(n1003), .ZN(n1005) );
  INV_X1 U1098 ( .A(G29), .ZN(n1004) );
  NAND2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1100 ( .A1(n1006), .A2(G11), .ZN(n1007) );
  XNOR2_X1 U1101 ( .A(n1007), .B(KEYINPUT121), .ZN(n1034) );
  XNOR2_X1 U1102 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1103 ( .A(n1008), .B(KEYINPUT122), .ZN(n1032) );
  XNOR2_X1 U1104 ( .A(n1009), .B(G1341), .ZN(n1014) );
  XOR2_X1 U1105 ( .A(G168), .B(G1966), .Z(n1010) );
  NOR2_X1 U1106 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1108 ( .A1(n1014), .A2(n1013), .ZN(n1030) );
  XNOR2_X1 U1109 ( .A(n1015), .B(KEYINPUT123), .ZN(n1017) );
  NAND2_X1 U1110 ( .A1(n1017), .A2(n1016), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(G171), .B(G1961), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(G303), .B(G1971), .ZN(n1019) );
  XNOR2_X1 U1113 ( .A(G299), .B(G1956), .ZN(n1018) );
  NOR2_X1 U1114 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1115 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XNOR2_X1 U1116 ( .A(G1348), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1117 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  NAND2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1120 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

