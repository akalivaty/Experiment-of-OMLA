//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n452), .A2(G567), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT65), .Z(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(new_n451), .B2(G2106), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n461), .A2(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(G162));
  OAI211_X1 g053(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n459), .A2(new_n460), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(KEYINPUT67), .ZN(new_n484));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n482), .A2(new_n486), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n481), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  XNOR2_X1  g069(.A(KEYINPUT5), .B(G543), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n495), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n495), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n498), .A2(new_n504), .ZN(G166));
  NAND3_X1  g080(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT7), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n508), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n500), .B(new_n502), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT70), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  AND2_X1   g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(new_n518), .B1(new_n495), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n522), .B2(KEYINPUT68), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT68), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n501), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(KEYINPUT69), .A3(G543), .A4(new_n524), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(G51), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n520), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND3_X1  g109(.A1(new_n526), .A2(G52), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n495), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n513), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G651), .B1(new_n540), .B2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n497), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n526), .A2(G43), .A3(new_n531), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n540), .A2(G81), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n546), .A2(KEYINPUT71), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT71), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n495), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n497), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(G91), .B2(new_n540), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n530), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n560));
  XNOR2_X1  g135(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n503), .B2(new_n527), .ZN(new_n564));
  NAND2_X1  g139(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n564), .A2(G53), .A3(new_n524), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n562), .A2(KEYINPUT73), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT73), .B1(new_n562), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND3_X1  g146(.A1(new_n564), .A2(G49), .A3(new_n524), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n495), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n540), .A2(G87), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n495), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n497), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n495), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n503), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G305));
  NAND3_X1  g157(.A1(new_n526), .A2(G47), .A3(new_n531), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n537), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n586), .A2(G651), .B1(new_n540), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT76), .B1(new_n513), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n526), .A2(G54), .A3(new_n531), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n495), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n497), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT77), .B1(new_n596), .B2(new_n598), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  XOR2_X1   g184(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n551), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n604), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT79), .Z(G323));
  XOR2_X1   g191(.A(G323), .B(KEYINPUT80), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n477), .A2(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n477), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n472), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT81), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT16), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT82), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n638), .A2(new_n640), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n638), .A2(new_n640), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT83), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(KEYINPUT83), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n653), .B(G14), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(KEYINPUT17), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n664), .B2(new_n661), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT87), .Z(new_n666));
  INV_X1    g241(.A(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n661), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n661), .A2(new_n660), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n666), .B(new_n670), .C1(new_n664), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G2096), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(G2096), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n622), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n672), .A2(G2096), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(G2100), .A3(new_n673), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n689), .A2(new_n691), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n687), .A2(new_n692), .A3(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT92), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n699), .B2(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n683), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n711), .A2(new_n682), .A3(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT23), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n608), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT107), .B(G1956), .Z(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT93), .B(G29), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G162), .B2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT29), .Z(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT106), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n720), .A2(G26), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT99), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n477), .A2(G140), .ZN(new_n733));
  NOR2_X1   g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT98), .Z(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n472), .A2(KEYINPUT97), .A3(G128), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT97), .B1(new_n472), .B2(G128), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n733), .B1(new_n735), .B2(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n732), .B1(G29), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT100), .B(G2067), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G33), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(new_n468), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT25), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G139), .B2(new_n477), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n744), .B1(new_n751), .B2(new_n743), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n720), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n470), .B2(new_n743), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2084), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n477), .A2(G141), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n472), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n743), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n743), .B2(G32), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n742), .A2(new_n753), .A3(new_n760), .A4(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n724), .A2(new_n725), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n721), .A2(G27), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n721), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n728), .A2(new_n771), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n714), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n551), .B2(new_n714), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n719), .B(new_n777), .C1(G1341), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G5), .A2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT103), .Z(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G301), .B2(new_n714), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n785), .B1(G2084), .B2(new_n759), .C1(new_n768), .C2(new_n769), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT105), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(new_n717), .B2(new_n718), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n780), .B(new_n788), .C1(new_n787), .C2(new_n786), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n779), .A2(G1341), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n714), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n604), .B2(new_n714), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n790), .B1(G1348), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G1348), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(G168), .A2(new_n714), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n714), .B2(G21), .ZN(new_n796));
  INV_X1    g371(.A(G1966), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT31), .B(G11), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n629), .A2(new_n720), .ZN(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n800), .B(new_n801), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n783), .A2(new_n784), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n796), .A2(new_n797), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n798), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT104), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n789), .A2(new_n794), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n714), .A2(G23), .ZN(new_n811));
  INV_X1    g386(.A(G288), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n714), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT33), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1976), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(G1976), .ZN(new_n817));
  INV_X1    g392(.A(G305), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n714), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G6), .B2(new_n714), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n714), .A2(G22), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G166), .B2(new_n714), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1971), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n816), .A2(new_n817), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n830));
  MUX2_X1   g405(.A(G24), .B(G290), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1986), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n477), .A2(G131), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n472), .A2(G119), .ZN(new_n835));
  NOR2_X1   g410(.A1(G95), .A2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT94), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n721), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G25), .B2(new_n721), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G1991), .Z(new_n842));
  OAI21_X1  g417(.A(new_n833), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g418(.A(new_n832), .B(new_n843), .C1(new_n842), .C2(new_n841), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n829), .A2(new_n830), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n810), .A2(new_n847), .A3(new_n848), .ZN(G311));
  NAND3_X1  g424(.A1(new_n810), .A2(new_n847), .A3(new_n848), .ZN(G150));
  NAND3_X1  g425(.A1(new_n526), .A2(G55), .A3(new_n531), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n537), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n854), .A2(G651), .B1(new_n540), .B2(G93), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n550), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n545), .B(new_n858), .C1(new_n548), .C2(new_n549), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT38), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n604), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n864), .A2(new_n865), .A3(G860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n856), .A2(G860), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n866), .A2(new_n868), .ZN(G145));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n629), .B(new_n470), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(G162), .Z(new_n872));
  XNOR2_X1  g447(.A(G164), .B(new_n739), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n766), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n766), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n750), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n751), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n477), .A2(G142), .ZN(new_n880));
  NOR2_X1   g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n472), .A2(KEYINPUT108), .A3(G130), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT108), .B1(new_n472), .B2(G130), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n880), .B1(new_n881), .B2(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n620), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n838), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n877), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n877), .B2(new_n879), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n872), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n872), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n870), .B(new_n892), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g474(.A(new_n614), .B(new_n860), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n603), .A2(new_n608), .ZN(new_n901));
  OAI211_X1 g476(.A(G299), .B(new_n595), .C1(new_n601), .C2(new_n602), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT41), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n900), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(KEYINPUT110), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(new_n818), .ZN(new_n911));
  NOR2_X1   g486(.A1(G290), .A2(G166), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G290), .A2(G166), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n910), .A2(new_n818), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n911), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n911), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n909), .B(new_n919), .ZN(new_n920));
  MUX2_X1   g495(.A(new_n856), .B(new_n920), .S(G868), .Z(G295));
  MUX2_X1   g496(.A(new_n856), .B(new_n920), .S(G868), .Z(G331));
  INV_X1    g497(.A(KEYINPUT114), .ZN(new_n923));
  INV_X1    g498(.A(new_n919), .ZN(new_n924));
  NOR2_X1   g499(.A1(G286), .A2(G301), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n520), .A2(new_n532), .B1(new_n535), .B2(new_n541), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n857), .A2(new_n859), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n857), .A2(KEYINPUT113), .A3(new_n927), .A4(new_n859), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n857), .B2(new_n859), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g510(.A(KEYINPUT112), .B(new_n927), .C1(new_n857), .C2(new_n859), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n932), .B(new_n903), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n928), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n905), .A2(new_n906), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n924), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n923), .B1(new_n940), .B2(G37), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n903), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT41), .ZN(new_n944));
  INV_X1    g519(.A(new_n927), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n546), .A2(new_n547), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT71), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n546), .A2(KEYINPUT71), .A3(new_n547), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n858), .B1(new_n950), .B2(new_n545), .ZN(new_n951));
  INV_X1    g526(.A(new_n859), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n943), .A2(new_n944), .B1(new_n953), .B2(new_n928), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n933), .A2(new_n934), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n955), .A2(new_n956), .B1(new_n930), .B2(new_n931), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n903), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT114), .B(new_n870), .C1(new_n958), .C2(new_n924), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n937), .A2(new_n924), .A3(new_n939), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n941), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n958), .B2(new_n924), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n956), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n907), .B1(new_n966), .B2(new_n932), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n953), .A2(new_n903), .A3(new_n928), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n919), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n965), .A3(new_n870), .A4(new_n960), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT115), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n963), .A2(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(KEYINPUT44), .C1(new_n961), .C2(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n461), .A2(new_n485), .A3(G2105), .ZN(new_n981));
  INV_X1    g556(.A(new_n489), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n487), .B(new_n492), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n479), .B(KEYINPUT66), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n464), .A2(new_n469), .A3(G40), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n739), .B(G2067), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT116), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n766), .B(G1996), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n842), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n838), .B(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n839), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n993), .A2(new_n994), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n739), .A2(G2067), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n988), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n991), .A2(new_n766), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n988), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n989), .A2(G1996), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT46), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(new_n1010), .C1(KEYINPUT46), .C2(new_n1008), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1005), .B1(KEYINPUT47), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1001), .B(new_n1013), .C1(KEYINPUT47), .C2(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT124), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G290), .B(G1986), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n997), .B1(new_n988), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n986), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n987), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n784), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n987), .B1(new_n985), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1024), .A2(KEYINPUT53), .A3(new_n775), .A4(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1022), .A2(KEYINPUT122), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT122), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT117), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1024), .A2(new_n1031), .A3(new_n1025), .ZN(new_n1032));
  AOI21_X1  g607(.A(G2078), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1027), .A2(new_n1028), .B1(new_n1033), .B2(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1032), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n775), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1022), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1026), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(G301), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT54), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n987), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n986), .A2(KEYINPUT121), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n985), .B2(new_n987), .ZN(new_n1049));
  AOI21_X1  g624(.A(G2067), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1348), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n603), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1956), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1021), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n562), .A2(new_n566), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n559), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1024), .A2(new_n1025), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1050), .A2(new_n1052), .A3(new_n603), .A4(KEYINPUT60), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT58), .B(G1341), .Z(new_n1070));
  NAND3_X1  g645(.A1(new_n1047), .A2(new_n1049), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1996), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1024), .A2(new_n1072), .A3(new_n1025), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n551), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1077), .A3(new_n551), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1069), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n604), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT60), .B1(new_n1054), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1068), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1045), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1034), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G301), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT54), .B(new_n1085), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n986), .B2(new_n1046), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n812), .A2(G1976), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT52), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n578), .A2(new_n681), .A3(new_n579), .A4(new_n581), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n580), .A2(new_n503), .ZN(new_n1102));
  OAI21_X1  g677(.A(G1981), .B1(new_n577), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT119), .B(KEYINPUT49), .C1(new_n1101), .C2(new_n1103), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1093), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1096), .B(new_n1099), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1971), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1030), .A2(new_n1111), .A3(new_n1032), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1019), .A2(new_n725), .A3(new_n1020), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT55), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n1118));
  NOR2_X1   g693(.A1(G166), .A2(new_n1092), .ZN(new_n1119));
  MUX2_X1   g694(.A(new_n1117), .B(new_n1118), .S(new_n1119), .Z(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1110), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1063), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1066), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1056), .A4(new_n1062), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1064), .A2(new_n1124), .A3(new_n1126), .A4(new_n1067), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n1092), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1029), .A2(new_n797), .ZN(new_n1131));
  INV_X1    g706(.A(G2084), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1019), .A2(new_n1132), .A3(new_n1020), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G168), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(G286), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1130), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1133), .A3(G168), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT51), .B1(new_n1138), .B2(G8), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1092), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1120), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1122), .A2(new_n1127), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1083), .A2(new_n1091), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1104), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1109), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1141), .B2(new_n1120), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1142), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1035), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1137), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1139), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT62), .A3(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n812), .A2(new_n1097), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1101), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1153), .A2(new_n1151), .B1(new_n1093), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1135), .A2(new_n1092), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1166), .A2(new_n1142), .A3(new_n1151), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1122), .A2(KEYINPUT63), .A3(new_n1142), .A4(new_n1167), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1145), .B(new_n1161), .C1(new_n1172), .C2(KEYINPUT120), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1164), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1015), .B(new_n1017), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  AND4_X1   g754(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1143), .A2(new_n1045), .A3(new_n1082), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1091), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1172), .A2(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1015), .B1(new_n1185), .B2(new_n1017), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1014), .B1(new_n1179), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g762(.A1(new_n676), .A2(new_n678), .A3(G319), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT126), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1191));
  NAND4_X1  g765(.A1(new_n676), .A2(new_n678), .A3(new_n1191), .A4(G319), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n1193), .A2(new_n710), .A3(new_n712), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n658), .A2(new_n1194), .A3(new_n898), .ZN(new_n1195));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n870), .B1(new_n958), .B2(new_n924), .ZN(new_n1197));
  AOI22_X1  g771(.A1(new_n1197), .A2(new_n923), .B1(new_n924), .B2(new_n958), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n965), .B1(new_n1198), .B2(new_n959), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n970), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1195), .B(new_n1196), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1196), .B1(new_n973), .B2(new_n1195), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  OAI21_X1  g778(.A(new_n1195), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1205), .A2(KEYINPUT127), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1206), .A2(new_n1201), .ZN(G225));
endmodule


