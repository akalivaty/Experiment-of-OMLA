//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(KEYINPUT3), .A3(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n477), .A2(new_n478), .A3(G137), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n468), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n478), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n479), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(G100), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(new_n479), .A3(KEYINPUT70), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT70), .B1(new_n488), .B2(new_n479), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n479), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND4_X1  g068(.A1(new_n477), .A2(new_n478), .A3(G126), .A4(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n479), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  AOI211_X1 g077(.A(new_n502), .B(new_n495), .C1(new_n497), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n494), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n477), .A2(new_n478), .A3(G138), .A4(new_n479), .ZN(new_n505));
  INV_X1    g080(.A(new_n465), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n507), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n505), .A2(KEYINPUT4), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT74), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n512), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT73), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(KEYINPUT6), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n517), .A2(new_n521), .A3(KEYINPUT75), .A4(new_n524), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n522), .A2(new_n523), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n535));
  AND2_X1   g110(.A1(KEYINPUT73), .A2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT73), .A2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT76), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n517), .A2(new_n521), .A3(G543), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n540), .A2(new_n542), .B1(G50), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n530), .A2(new_n544), .ZN(G303));
  INV_X1    g120(.A(G303), .ZN(G166));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(G89), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n527), .A2(new_n528), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G63), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n522), .B2(new_n523), .ZN(new_n550));
  AND3_X1   g125(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n517), .A2(new_n521), .A3(G51), .A4(G543), .ZN(new_n553));
  NAND3_X1  g128(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n548), .A2(new_n557), .ZN(G168));
  NAND3_X1  g133(.A1(new_n527), .A2(G90), .A3(new_n528), .ZN(new_n559));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n522), .B2(new_n523), .ZN(new_n561));
  AND2_X1   g136(.A1(G77), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n539), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(G52), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n517), .A2(new_n521), .A3(G543), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n559), .A2(new_n566), .ZN(G171));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n522), .B2(new_n523), .ZN(new_n569));
  AND2_X1   g144(.A1(G68), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n539), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT79), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n539), .B(new_n573), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n527), .A2(G81), .A3(new_n528), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(G43), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n543), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT81), .ZN(G176));
  NAND2_X1  g157(.A1(G1), .A2(G3), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT8), .ZN(new_n584));
  NAND4_X1  g159(.A1(G319), .A2(G483), .A3(G661), .A4(new_n584), .ZN(G188));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT83), .B(G65), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n527), .A2(G91), .A3(new_n528), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n538), .A2(KEYINPUT6), .B1(new_n513), .B2(new_n516), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n591), .A2(new_n592), .A3(G53), .A4(G543), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n517), .A2(new_n521), .A3(G53), .A4(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n593), .A2(KEYINPUT82), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT82), .B1(new_n593), .B2(new_n595), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n589), .B(new_n590), .C1(new_n596), .C2(new_n597), .ZN(G299));
  NAND2_X1  g173(.A1(new_n559), .A2(new_n566), .ZN(G301));
  NAND2_X1  g174(.A1(new_n548), .A2(new_n557), .ZN(G286));
  NAND3_X1  g175(.A1(new_n527), .A2(G87), .A3(new_n528), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n524), .A2(G74), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n543), .A2(G49), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(G288));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n532), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n543), .A2(G48), .B1(new_n607), .B2(new_n539), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n527), .A2(G86), .A3(new_n528), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n543), .A2(G47), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n527), .A2(new_n528), .ZN(new_n613));
  INV_X1    g188(.A(G85), .ZN(new_n614));
  OAI221_X1 g189(.A(new_n611), .B1(new_n538), .B2(new_n612), .C1(new_n613), .C2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n527), .A2(G92), .A3(new_n528), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n527), .A2(new_n619), .A3(G92), .A4(new_n528), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n532), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n543), .A2(G54), .B1(new_n623), .B2(G651), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n616), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G299), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  XNOR2_X1  g205(.A(G280), .B(KEYINPUT84), .ZN(G297));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND3_X1  g208(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(G559), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n484), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n486), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n479), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n506), .A2(new_n472), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT13), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n689), .B(new_n688), .S(new_n681), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(G301), .A2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G5), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G1961), .ZN(new_n703));
  NAND2_X1  g278(.A1(G160), .A2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n705), .B2(KEYINPUT24), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(KEYINPUT24), .B2(new_n705), .ZN(new_n707));
  AOI21_X1  g282(.A(G2084), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G32), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G141), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n472), .A2(G105), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G129), .B2(new_n486), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n710), .B1(new_n720), .B2(new_n709), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  AOI211_X1 g297(.A(new_n703), .B(new_n708), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n709), .A2(G33), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n506), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(new_n479), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n484), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n709), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G2072), .Z(new_n734));
  NAND3_X1  g309(.A1(new_n704), .A2(G2084), .A3(new_n707), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(new_n721), .C2(new_n722), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT93), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n709), .A2(G35), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT95), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n709), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT97), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g321(.A1(new_n724), .A2(new_n737), .A3(new_n738), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT98), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n709), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n709), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G28), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n709), .B1(new_n756), .B2(G28), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n755), .B1(new_n757), .B2(new_n758), .C1(new_n645), .C2(new_n709), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n699), .A2(G21), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G286), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n701), .A2(new_n760), .B1(new_n763), .B2(G1966), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n709), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n486), .A2(G128), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n479), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OR4_X1    g349(.A1(new_n754), .A2(new_n759), .A3(new_n764), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n625), .A2(new_n699), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G4), .B2(new_n699), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n699), .A2(G19), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n579), .B2(new_n699), .ZN(new_n781));
  AOI22_X1  g356(.A1(G1341), .A2(new_n781), .B1(new_n763), .B2(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n777), .A2(new_n778), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n782), .B(new_n783), .C1(G1341), .C2(new_n781), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n751), .A2(new_n775), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n699), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n629), .B2(new_n699), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT99), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n747), .A2(new_n750), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(KEYINPUT91), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(G290), .B(KEYINPUT88), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G16), .B2(G24), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT89), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT89), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G1986), .ZN(new_n801));
  NOR2_X1   g376(.A1(G25), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n484), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n486), .A2(G119), .ZN(new_n804));
  OR2_X1    g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT87), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  INV_X1    g387(.A(G1986), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n798), .B2(new_n799), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n801), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n699), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n699), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1971), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n699), .A2(G23), .ZN(new_n819));
  INV_X1    g394(.A(G288), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n699), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT33), .B(G1976), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT90), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G6), .A2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G305), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT32), .B(G1981), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n818), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  AOI21_X1  g406(.A(new_n794), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n815), .A2(new_n794), .A3(new_n831), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n791), .B1(new_n833), .B2(new_n834), .ZN(G311));
  INV_X1    g410(.A(new_n791), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n832), .ZN(G150));
  NOR2_X1   g413(.A1(new_n634), .A2(new_n632), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n527), .A2(G93), .A3(new_n528), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n543), .A2(G55), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n532), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n539), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT101), .B1(new_n849), .B2(new_n539), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n842), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n856), .A2(new_n579), .A3(new_n846), .A4(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n841), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT104), .ZN(G145));
  XNOR2_X1  g442(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n510), .B(new_n771), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n720), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n720), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n732), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n731), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n484), .A2(G142), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n486), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n479), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n648), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n808), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n645), .B(G160), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n492), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n874), .A2(new_n876), .A3(new_n889), .A4(new_n884), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n874), .A2(new_n876), .A3(new_n884), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT106), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n884), .B1(new_n874), .B2(new_n876), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n888), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n869), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n892), .ZN(new_n901));
  INV_X1    g476(.A(new_n888), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n894), .A3(new_n868), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n904), .ZN(G395));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n858), .B(new_n636), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n625), .A2(G299), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT82), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT82), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n590), .A2(new_n589), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n634), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n908), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n625), .A2(G299), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n908), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n906), .B1(new_n907), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n858), .B(new_n635), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(KEYINPUT109), .A3(new_n921), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n918), .A2(new_n920), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n907), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  XNOR2_X1  g507(.A(G288), .B(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G303), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  XNOR2_X1  g510(.A(G288), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G166), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G290), .B(G305), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n938), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n925), .A2(new_n927), .A3(new_n942), .A4(new_n930), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n932), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n932), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n853), .A2(new_n854), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(G868), .B2(new_n947), .ZN(G295));
  OAI21_X1  g523(.A(new_n946), .B1(G868), .B2(new_n947), .ZN(G331));
  AOI21_X1  g524(.A(G286), .B1(G171), .B2(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(G301), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT111), .B(KEYINPUT112), .C1(new_n559), .C2(new_n566), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n559), .A2(KEYINPUT111), .A3(new_n566), .ZN(new_n956));
  NAND2_X1  g531(.A1(G168), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G301), .A2(new_n952), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT112), .ZN(new_n959));
  NAND3_X1  g534(.A1(G301), .A2(new_n952), .A3(new_n951), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n858), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(G168), .B(new_n956), .C1(new_n953), .C2(new_n954), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n957), .A3(new_n960), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n855), .A4(new_n857), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n921), .A2(new_n923), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n962), .A2(new_n928), .A3(new_n965), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n941), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n962), .A2(new_n965), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n924), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n938), .A2(new_n940), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n939), .B1(new_n934), .B2(new_n937), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n962), .A2(new_n928), .A3(new_n965), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  INV_X1    g553(.A(G37), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n908), .A2(new_n917), .ZN(new_n984));
  AND4_X1   g559(.A1(new_n855), .A2(new_n963), .A3(new_n964), .A4(new_n857), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n963), .A2(new_n964), .B1(new_n855), .B2(new_n857), .ZN(new_n986));
  OAI211_X1 g561(.A(KEYINPUT41), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n922), .B1(new_n962), .B2(new_n965), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(new_n975), .C1(new_n929), .C2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n968), .A3(new_n979), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n990), .B2(KEYINPUT43), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n982), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT114), .B1(new_n982), .B2(new_n991), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n968), .B1(new_n980), .B2(new_n981), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(KEYINPUT43), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n992), .A2(new_n993), .B1(new_n996), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g572(.A(new_n807), .B(new_n810), .Z(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT115), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n771), .B(new_n773), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n720), .A2(G1996), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n719), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(G290), .B(new_n813), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n504), .B2(new_n509), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n468), .A2(G40), .A3(new_n473), .A4(new_n480), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  INV_X1    g590(.A(G1966), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1010), .A2(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n504), .B2(new_n509), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1012), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1012), .B1(new_n510), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2084), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1015), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT118), .B(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G168), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT51), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(KEYINPUT51), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(KEYINPUT125), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1029), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(KEYINPUT125), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1030), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n601), .A2(new_n603), .A3(G1976), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1036), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n820), .B2(G1976), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G305), .A2(G1981), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n608), .B2(new_n609), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT119), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n1048), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1049), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n510), .A2(new_n1008), .A3(new_n1020), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1036), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1047), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1019), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT116), .B(new_n1018), .C1(new_n504), .C2(new_n509), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1011), .A2(new_n1063), .A3(new_n1020), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT117), .B(G1971), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1024), .A2(new_n745), .A3(new_n1026), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1061), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1069), .B2(new_n1036), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1065), .B2(G2078), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1078));
  INV_X1    g653(.A(G2078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n760), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1074), .A2(new_n1075), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT127), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1041), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1041), .B2(new_n1085), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1039), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G288), .A2(G1976), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1049), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1061), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1093), .A2(new_n1059), .B1(new_n1094), .B2(new_n1073), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n1096), .B2(new_n1015), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1072), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1069), .A2(new_n1099), .A3(G8), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1074), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1033), .A2(G168), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1103), .A2(KEYINPUT63), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1098), .B1(new_n1096), .B2(new_n1029), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(new_n1103), .A3(new_n1073), .A4(new_n1061), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1095), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1011), .A2(new_n1063), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1020), .A3(new_n1064), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n910), .A2(new_n911), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n915), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT122), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n914), .A2(KEYINPUT57), .A3(new_n916), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n1115), .C1(new_n915), .C2(new_n1116), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1956), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AND4_X1   g699(.A1(new_n1111), .A2(new_n1114), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1114), .A2(new_n1124), .A3(new_n1122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1348), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1009), .A2(G2067), .A3(new_n1012), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n625), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1122), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1113), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1065), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(new_n1123), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1126), .A2(new_n1128), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1058), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1065), .B2(G1996), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n579), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n579), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1130), .B1(new_n1081), .B2(new_n778), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n634), .B1(new_n1146), .B2(KEYINPUT60), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  NOR4_X1   g723(.A1(new_n1129), .A2(new_n1148), .A3(new_n625), .A4(new_n1130), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1147), .A2(new_n1149), .B1(KEYINPUT60), .B2(new_n1146), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1135), .A2(new_n1127), .A3(KEYINPUT61), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1145), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1134), .A2(new_n1123), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1111), .B1(new_n1153), .B2(new_n1122), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1135), .B1(new_n1154), .B2(new_n1125), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1136), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G301), .B(KEYINPUT54), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1112), .A2(new_n1064), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1079), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n480), .A2(new_n473), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n467), .A2(KEYINPUT126), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n479), .B1(new_n467), .B2(KEYINPUT126), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1163), .B(new_n1164), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1161), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1160), .A2(new_n1168), .B1(new_n1083), .B2(new_n1161), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1159), .A2(new_n1106), .A3(new_n1102), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1110), .B1(new_n1158), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1014), .B1(new_n1090), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1000), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1013), .B1(new_n1173), .B2(new_n719), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1013), .A2(new_n1002), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1175), .A2(KEYINPUT46), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(KEYINPUT46), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT47), .Z(new_n1179));
  INV_X1    g754(.A(new_n1013), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1180), .A2(G1986), .A3(G290), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1005), .A2(new_n1180), .B1(KEYINPUT48), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(KEYINPUT48), .B2(new_n1181), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n808), .A2(new_n810), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1004), .A2(new_n1184), .B1(G2067), .B2(new_n771), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1179), .B(new_n1183), .C1(new_n1013), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g762(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G229), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g764(.A(new_n1190), .B1(new_n895), .B2(new_n899), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1191), .A2(new_n996), .ZN(G308));
  NAND2_X1  g766(.A1(new_n903), .A2(new_n894), .ZN(new_n1193));
  AND2_X1   g767(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n1193), .B(new_n1190), .C1(new_n1194), .C2(new_n994), .ZN(G225));
endmodule


