//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n469), .A2(new_n466), .A3(G101), .A4(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(G137), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(new_n482));
  AOI21_X1  g057(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n480), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n466), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n463), .A2(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G138), .A4(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n483), .A2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n466), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT70), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  AOI211_X1 g077(.A(new_n502), .B(new_n499), .C1(new_n494), .C2(new_n497), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n492), .B(new_n493), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n512), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT73), .Z(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n508), .A2(new_n531), .B1(new_n510), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n514), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n508), .A2(new_n537), .B1(new_n510), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n514), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  AND2_X1   g125(.A1(KEYINPUT6), .A2(G651), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT6), .A2(G651), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n559), .A2(new_n514), .B1(new_n508), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  AND2_X1   g141(.A1(G49), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n507), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n551), .C2(new_n552), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(G74), .A2(G651), .ZN(new_n573));
  AND2_X1   g148(.A1(KEYINPUT5), .A2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT5), .A2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n514), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT76), .B(G651), .C1(new_n506), .C2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n506), .A2(new_n507), .A3(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n571), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n508), .A2(new_n582), .B1(new_n510), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n514), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n508), .A2(new_n589), .B1(new_n510), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n514), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n591), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n506), .A2(new_n507), .A3(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT10), .Z(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n598), .A2(new_n554), .A3(KEYINPUT77), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT77), .B1(new_n598), .B2(new_n554), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n576), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n555), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n595), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n595), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n562), .ZN(G280));
  XNOR2_X1  g184(.A(G280), .B(KEYINPUT78), .ZN(G297));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n605), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n605), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n545), .B2(G868), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n465), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n483), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n466), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT79), .B(G2100), .Z(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n640), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n651), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n648), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n666), .A2(KEYINPUT20), .A3(new_n670), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n671), .B1(new_n670), .B2(new_n667), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G35), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G162), .B2(G29), .ZN(new_n686));
  INV_X1    g261(.A(G2090), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G26), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(G116), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G2105), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT94), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n483), .A2(G128), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n465), .A2(G140), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n693), .B1(new_n701), .B2(new_n691), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2067), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n691), .A2(G32), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT96), .Z(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(KEYINPUT26), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(KEYINPUT26), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n483), .A2(G129), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n465), .A2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n704), .B1(new_n713), .B2(new_n691), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT27), .B(G1996), .Z(new_n715));
  AOI21_X1  g290(.A(new_n703), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G4), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n605), .B2(G16), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n690), .B(new_n716), .C1(G1348), .C2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n545), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(G19), .ZN(new_n722));
  INV_X1    g297(.A(G1341), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n720), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n722), .A2(new_n723), .B1(G1966), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n720), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n720), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G34), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n476), .B2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n718), .A2(G1348), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR2_X1   g316(.A1(new_n621), .A2(new_n691), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT30), .B(G28), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n741), .B(new_n742), .C1(new_n691), .C2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n726), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n691), .A2(G33), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n489), .A2(G127), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n466), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n749), .B(new_n752), .C1(G139), .C2(new_n465), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT95), .Z(new_n754));
  AOI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n722), .A2(new_n723), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n691), .A2(G27), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n504), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT99), .B(G2078), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n725), .A2(G1966), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n746), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n714), .A2(new_n715), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT97), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n688), .B2(new_n689), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n720), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n562), .B2(new_n720), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1956), .Z(new_n770));
  OAI221_X1 g345(.A(new_n770), .B1(new_n760), .B2(new_n761), .C1(new_n756), .C2(new_n755), .ZN(new_n771));
  OR4_X1    g346(.A1(new_n719), .A2(new_n763), .A3(new_n766), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n720), .A2(G23), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n577), .A2(new_n578), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n580), .B1(new_n568), .B2(new_n570), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n571), .A2(new_n579), .A3(KEYINPUT92), .A4(new_n580), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(new_n720), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n720), .A2(G22), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n720), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G1971), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(G1971), .ZN(new_n787));
  NOR2_X1   g362(.A1(G6), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n587), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n789), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n691), .A2(G25), .ZN(new_n797));
  OR2_X1    g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT87), .ZN(new_n800));
  AOI22_X1  g375(.A1(G119), .A2(new_n483), .B1(new_n465), .B2(G131), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n691), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT88), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(KEYINPUT89), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(KEYINPUT89), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n720), .A2(G24), .ZN(new_n810));
  INV_X1    g385(.A(G290), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n720), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n795), .A2(new_n796), .A3(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT36), .Z(new_n816));
  NOR2_X1   g391(.A1(new_n772), .A2(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  NAND2_X1  g393(.A1(new_n605), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT103), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n506), .A2(new_n507), .A3(G93), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT101), .B(G55), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n822), .B1(new_n510), .B2(new_n823), .C1(new_n824), .C2(new_n514), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n541), .B2(new_n539), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n543), .A2(new_n544), .A3(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n821), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  INV_X1    g408(.A(new_n826), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(G145));
  XOR2_X1   g412(.A(new_n701), .B(new_n504), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n713), .ZN(new_n839));
  MUX2_X1   g414(.A(new_n753), .B(new_n754), .S(new_n839), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n802), .B(new_n624), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n483), .A2(G130), .ZN(new_n842));
  OR2_X1    g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n465), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n841), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n840), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n621), .B(new_n476), .ZN(new_n851));
  XOR2_X1   g426(.A(G162), .B(new_n851), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  INV_X1    g429(.A(new_n852), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n848), .A2(new_n855), .A3(new_n849), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n562), .A2(new_n604), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT104), .ZN(new_n861));
  NAND2_X1  g436(.A1(G299), .A2(new_n605), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n859), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n860), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n829), .B(new_n613), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT105), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n866), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n862), .A2(new_n860), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n779), .B(new_n587), .ZN(new_n878));
  XNOR2_X1  g453(.A(G166), .B(new_n811), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n870), .A2(new_n881), .A3(new_n873), .A4(new_n875), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n877), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(G868), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n826), .A2(G868), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(G295));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(G331));
  INV_X1    g463(.A(new_n880), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT106), .B1(new_n874), .B2(new_n859), .ZN(new_n890));
  INV_X1    g465(.A(new_n861), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n865), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n874), .A2(KEYINPUT106), .A3(new_n859), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n827), .A2(new_n828), .A3(G301), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G301), .B1(new_n827), .B2(new_n828), .ZN(new_n896));
  OAI21_X1  g471(.A(G286), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(G168), .A3(new_n894), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n892), .A2(new_n893), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n897), .A2(new_n899), .A3(new_n874), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n889), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n899), .A3(new_n874), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n897), .A2(new_n899), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n880), .B(new_n903), .C1(new_n904), .C2(new_n867), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .A4(new_n854), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n899), .A2(new_n897), .B1(new_n864), .B2(new_n866), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n880), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n906), .A4(new_n902), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(new_n880), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n905), .A2(new_n854), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n906), .B1(new_n914), .B2(new_n915), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n902), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n493), .B1(new_n501), .B2(new_n503), .ZN(new_n926));
  INV_X1    g501(.A(new_n492), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n471), .A2(new_n475), .A3(G40), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT108), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n471), .A2(new_n475), .A3(new_n933), .A4(G40), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G2067), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n701), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT109), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n713), .B(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n803), .A2(new_n805), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n803), .A2(new_n805), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G1986), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n936), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n932), .A2(new_n504), .A3(new_n925), .A4(new_n934), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n947), .A2(G8), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT112), .A4(G1976), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n777), .A2(new_n778), .A3(G1976), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1976), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(G288), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n948), .A2(new_n949), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1981), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n587), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n584), .A2(new_n586), .A3(G1981), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(KEYINPUT49), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n957), .B2(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n948), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n948), .A2(KEYINPUT113), .A3(new_n952), .A4(new_n949), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n932), .A2(new_n934), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n930), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT110), .B(G1971), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n504), .B2(new_n925), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(new_n935), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n504), .A2(new_n978), .A3(new_n925), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n687), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n972), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n517), .A2(G8), .A3(new_n518), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT55), .Z(new_n985));
  OR2_X1    g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n983), .A2(new_n987), .A3(new_n985), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n983), .B2(new_n985), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n971), .B(new_n986), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n928), .A2(KEYINPUT50), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n973), .A3(new_n981), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n992), .A2(KEYINPUT115), .B1(new_n995), .B2(new_n731), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n975), .A2(new_n997), .A3(new_n991), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(G8), .A3(G168), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n946), .B1(new_n990), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n971), .A2(new_n986), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n983), .A2(new_n985), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n972), .B(G286), .C1(new_n996), .C2(new_n998), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1002), .A2(KEYINPUT116), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1001), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n988), .A2(new_n989), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1011), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n971), .A2(new_n986), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(KEYINPUT117), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(KEYINPUT117), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n996), .A2(G168), .A3(new_n998), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT51), .ZN(new_n1020));
  AOI21_X1  g595(.A(G168), .B1(new_n996), .B2(new_n998), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n1018), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT62), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2078), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n930), .A2(new_n973), .A3(new_n1028), .A4(new_n974), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n994), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n993), .A2(new_n973), .A3(KEYINPUT118), .A4(new_n981), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n729), .A3(new_n1034), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1031), .B1(new_n1037), .B2(KEYINPUT123), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  AOI21_X1  g615(.A(G301), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n990), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1025), .A2(new_n1027), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G288), .A2(G1976), .ZN(new_n1044));
  XOR2_X1   g619(.A(new_n1044), .B(KEYINPUT114), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n964), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n960), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1011), .A2(new_n971), .B1(new_n948), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1017), .A2(new_n1043), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n990), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n930), .A2(new_n974), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT124), .B(G2078), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n931), .A2(new_n1030), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1052), .A2(new_n1054), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1035), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1041), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1038), .A2(G301), .A3(new_n1040), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1059), .B(new_n1062), .C1(new_n1061), .C2(new_n1060), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1050), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1348), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1033), .A2(new_n1065), .A3(new_n1034), .ZN(new_n1066));
  INV_X1    g641(.A(new_n947), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n937), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(KEYINPUT60), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n605), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1072), .A3(new_n605), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT60), .A4(new_n604), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n1069), .B2(new_n605), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1074), .A2(new_n1079), .B1(KEYINPUT60), .B2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n562), .A2(KEYINPUT57), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n558), .B2(new_n561), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1956), .B1(new_n980), .B2(new_n981), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  AND4_X1   g662(.A1(new_n973), .A2(new_n930), .A3(new_n974), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n930), .A2(new_n973), .A3(new_n974), .A4(new_n1087), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1084), .B(new_n1090), .C1(new_n995), .C2(G1956), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1091), .A3(KEYINPUT61), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .A4(KEYINPUT61), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT58), .B(G1341), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n975), .A2(G1996), .B1(new_n1067), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n545), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1103), .A3(new_n545), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1097), .A2(new_n1098), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1096), .A2(new_n1108), .A3(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1080), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1089), .B1(new_n1075), .B2(new_n604), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1091), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1064), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n945), .B1(new_n1049), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n936), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT48), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G290), .A2(G1986), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT48), .B1(new_n936), .B2(new_n1117), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1119), .B(new_n1120), .C1(new_n943), .C2(new_n936), .ZN(new_n1121));
  INV_X1    g696(.A(G1996), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT46), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n939), .A2(new_n713), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT46), .B1(new_n936), .B2(new_n1122), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1124), .A2(new_n1115), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT47), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n701), .A2(new_n937), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n939), .A2(new_n940), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n941), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1121), .B(new_n1129), .C1(new_n936), .C2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1114), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(G319), .ZN(new_n1136));
  NOR4_X1   g710(.A1(G229), .A2(new_n1136), .A3(G401), .A4(G227), .ZN(new_n1137));
  NAND3_X1  g711(.A1(new_n917), .A2(new_n1137), .A3(new_n857), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


