//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT69), .B(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n463), .B2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n464), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  AND4_X1   g051(.A1(G137), .A2(new_n474), .A3(new_n471), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n482), .B2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G125), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n478), .A2(new_n490), .ZN(G160));
  NAND2_X1  g066(.A1(new_n474), .A2(new_n476), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT71), .Z(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(new_n471), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G124), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(G162));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n474), .A2(new_n476), .A3(new_n502), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(KEYINPUT4), .B1(new_n481), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n474), .A2(G126), .A3(G2105), .A4(new_n476), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(G62), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n516), .A2(new_n517), .B1(new_n520), .B2(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n513), .A2(new_n512), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(new_n519), .A3(KEYINPUT72), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(G88), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n518), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G166));
  AND3_X1   g106(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AOI211_X1 g109(.A(new_n532), .B(new_n534), .C1(G51), .C2(new_n520), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(new_n528), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  XOR2_X1   g115(.A(KEYINPUT74), .B(G52), .Z(new_n541));
  NAND2_X1  g116(.A1(new_n520), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n542), .B1(new_n511), .B2(new_n543), .C1(new_n536), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n537), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n512), .A2(new_n513), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT76), .B(G43), .ZN(new_n553));
  AOI22_X1  g128(.A1(G651), .A2(new_n552), .B1(new_n520), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n526), .A2(G91), .A3(new_n528), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n520), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n519), .A2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT77), .B(new_n563), .C1(new_n569), .C2(new_n565), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n550), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n562), .A2(new_n568), .A3(new_n570), .A4(new_n574), .ZN(G299));
  XNOR2_X1  g150(.A(new_n545), .B(KEYINPUT75), .ZN(G301));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n530), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n518), .A2(new_n521), .A3(KEYINPUT78), .A4(new_n529), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G303));
  NAND3_X1  g155(.A1(new_n526), .A2(G87), .A3(new_n528), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n526), .A2(KEYINPUT79), .A3(G87), .A4(new_n528), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n527), .A2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n586), .A2(new_n511), .B1(new_n569), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n526), .A2(G86), .A3(new_n528), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G61), .B1(new_n512), .B2(new_n513), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT80), .B1(new_n596), .B2(G651), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n598), .B(new_n511), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n595), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n527), .B2(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n598), .B1(new_n602), .B2(new_n511), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n596), .A2(KEYINPUT80), .A3(G651), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n593), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n520), .A2(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(G85), .ZN(new_n611));
  OAI221_X1 g186(.A(new_n609), .B1(new_n511), .B2(new_n610), .C1(new_n536), .C2(new_n611), .ZN(G290));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G301), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n526), .A2(G92), .A3(new_n528), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n550), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(G651), .A2(new_n620), .B1(new_n520), .B2(G54), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n621), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n614), .B1(new_n613), .B2(new_n626), .ZN(G284));
  AOI21_X1  g202(.A(new_n614), .B1(new_n613), .B2(new_n626), .ZN(G321));
  NAND2_X1  g203(.A1(G299), .A2(new_n613), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G168), .B2(new_n613), .ZN(G280));
  XOR2_X1   g205(.A(G280), .B(KEYINPUT84), .Z(G297));
  XOR2_X1   g206(.A(KEYINPUT85), .B(G559), .Z(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(G860), .B2(new_n632), .ZN(G148));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n464), .A2(new_n472), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n481), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n493), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n498), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n471), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  INV_X1    g247(.A(new_n669), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n673), .B2(new_n667), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n667), .B(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n674), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n673), .A3(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G19), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n556), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1341), .Z(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G26), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  AND2_X1   g280(.A1(new_n474), .A2(new_n476), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(G140), .A3(new_n471), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n493), .A2(new_n709), .A3(G140), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(G128), .A3(G2105), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n705), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT91), .B(G2067), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n703), .A2(G27), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT99), .Z(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n703), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n702), .B(new_n720), .C1(G2078), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n703), .A2(G33), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n493), .A2(G139), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n729), .C1(new_n471), .C2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n703), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n699), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT23), .ZN(new_n737));
  INV_X1    g312(.A(G299), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n699), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G5), .A2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT97), .Z(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G301), .B2(new_n699), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n718), .B2(new_n719), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n733), .A2(G2072), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n724), .A2(new_n742), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n699), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n626), .B2(new_n699), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n699), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n699), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1966), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n745), .A2(new_n746), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n703), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n649), .B2(new_n703), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n758), .A2(new_n759), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT98), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n703), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n703), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT29), .B(G2090), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G160), .B2(new_n703), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT94), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2084), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n493), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n498), .A2(G129), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n638), .A2(G105), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT26), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(new_n703), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n703), .B2(G32), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT95), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n787), .A2(new_n789), .B1(G2078), .B2(new_n723), .ZN(new_n791));
  AND4_X1   g366(.A1(new_n771), .A2(new_n778), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n755), .A2(new_n767), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n493), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n498), .A2(G119), .ZN(new_n795));
  OR2_X1    g370(.A1(G95), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G25), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT35), .B(G1991), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n804), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n699), .A2(G24), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G290), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G1986), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n805), .A2(new_n806), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(G305), .A2(G16), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n699), .A2(G6), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT32), .B(G1981), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n817), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT89), .B1(new_n585), .B2(new_n589), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n825), .B(new_n588), .C1(new_n583), .C2(new_n584), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G16), .B2(G23), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT33), .B(G1976), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n699), .A2(G22), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G166), .B2(new_n699), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1971), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n829), .B2(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n823), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n812), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT34), .B1(new_n836), .B2(new_n823), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n793), .B1(new_n842), .B2(new_n844), .ZN(G311));
  INV_X1    g420(.A(G311), .ZN(G150));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n550), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(G651), .A2(new_n849), .B1(new_n520), .B2(G55), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(new_n536), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n555), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n555), .A2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n626), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT102), .ZN(new_n862));
  AOI21_X1  g437(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n853), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n493), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n498), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n471), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n640), .B(new_n873), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n717), .A2(G164), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n715), .B1(new_n708), .B2(new_n710), .ZN(new_n877));
  INV_X1    g452(.A(G164), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n876), .A2(new_n785), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n785), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n732), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n879), .ZN(new_n883));
  INV_X1    g458(.A(new_n785), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n876), .A2(new_n785), .A3(new_n879), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n731), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n887), .A3(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n885), .A2(new_n889), .A3(new_n731), .A4(new_n886), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n888), .A2(new_n798), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n798), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n875), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n799), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n798), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n874), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(G160), .B(new_n649), .Z(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(G162), .Z(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n893), .B2(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(KEYINPUT40), .A3(new_n901), .A4(new_n900), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(G395));
  XOR2_X1   g482(.A(new_n634), .B(new_n856), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n622), .B(new_n738), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT41), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n827), .B(G290), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n607), .B(G166), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT104), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n908), .A2(new_n910), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n920), .B(new_n921), .C1(new_n909), .C2(new_n908), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n913), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n919), .B1(new_n913), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n853), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n926), .ZN(G295));
  OAI21_X1  g502(.A(new_n925), .B1(G868), .B2(new_n926), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(G286), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G168), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n856), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n854), .A4(new_n855), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n935), .B2(new_n910), .ZN(new_n936));
  INV_X1    g511(.A(new_n909), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n918), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n936), .A2(new_n917), .A3(new_n916), .A4(new_n938), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n929), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n929), .A3(new_n941), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n940), .A2(new_n929), .A3(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(G397));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n505), .B2(new_n509), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n638), .A2(G101), .ZN(new_n955));
  INV_X1    g530(.A(new_n477), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n490), .A2(G40), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n884), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT107), .Z(new_n962));
  XNOR2_X1  g537(.A(new_n877), .B(G2067), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n959), .B2(new_n785), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n799), .A2(new_n804), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n798), .A2(new_n803), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n958), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(G1986), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n958), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n478), .A2(G40), .A3(new_n490), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n951), .C1(new_n505), .C2(new_n509), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n954), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT108), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n980));
  NOR2_X1   g555(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n505), .B2(new_n509), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(G40), .A3(new_n478), .A4(new_n490), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT109), .B(G2090), .Z(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT110), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n972), .A2(new_n987), .A3(new_n982), .A4(new_n985), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n977), .A2(new_n979), .A3(new_n986), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n578), .A2(G8), .A3(new_n579), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n578), .A2(KEYINPUT55), .A3(G8), .A4(new_n579), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT111), .B(G86), .Z(new_n1000));
  NAND3_X1  g575(.A1(new_n526), .A2(new_n528), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT112), .B1(new_n1001), .B2(new_n592), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n603), .A2(new_n604), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(KEYINPUT112), .A3(new_n592), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n999), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(G1981), .B(new_n593), .C1(new_n600), .C2(new_n606), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n607), .A2(new_n999), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1005), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1010), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1009), .B(KEYINPUT49), .C1(new_n1011), .C2(new_n999), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n957), .B2(new_n952), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n824), .A2(new_n826), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1013), .ZN(new_n1018));
  INV_X1    g593(.A(new_n824), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n585), .A2(KEYINPUT89), .A3(new_n589), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(G1976), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1016), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1014), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1015), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n995), .A2(new_n996), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n991), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G168), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n983), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n987), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n974), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n972), .A2(new_n987), .A3(new_n982), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT114), .B1(new_n1038), .B2(G2084), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1029), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n997), .A2(new_n1026), .A3(new_n1028), .A4(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1015), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n976), .A2(new_n988), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1027), .B1(new_n1043), .B2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1028), .A2(new_n1042), .A3(new_n1045), .A4(new_n1040), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1025), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1041), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  AND4_X1   g626(.A1(new_n1051), .A2(new_n1028), .A3(new_n1042), .A4(new_n1045), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1024), .A2(new_n1044), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT58), .B(G1341), .Z(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n957), .B2(new_n952), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(G1996), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n972), .A2(new_n954), .A3(new_n973), .A4(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT119), .B(new_n1056), .C1(new_n957), .C2(new_n952), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n556), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n556), .A3(new_n1065), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1038), .A2(new_n753), .ZN(new_n1070));
  INV_X1    g645(.A(G2067), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n972), .A2(new_n951), .A3(new_n1071), .A4(new_n878), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n626), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n626), .A2(KEYINPUT60), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1038), .A2(new_n740), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NAND3_X1  g657(.A1(G299), .A2(new_n1082), .A3(KEYINPUT57), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(G299), .B2(new_n1082), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n972), .A2(new_n954), .A3(new_n973), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1081), .A2(new_n1088), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n1084), .A2(KEYINPUT117), .A3(new_n1085), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT117), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT61), .B(new_n1089), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1089), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1086), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1069), .A2(new_n1080), .A3(new_n1094), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1076), .A2(new_n626), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1089), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT122), .B(new_n746), .C1(new_n980), .C2(new_n983), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT122), .B1(new_n1038), .B2(new_n746), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G2078), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n972), .A2(new_n954), .A3(new_n1108), .A4(new_n973), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(G2078), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G40), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n487), .B2(G2105), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n954), .A2(new_n478), .A3(new_n973), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1107), .A2(G301), .A3(new_n1112), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n746), .B1(new_n980), .B2(new_n983), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n972), .A2(new_n954), .A3(new_n973), .A4(new_n1113), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G171), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT121), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(G171), .C1(new_n1111), .C2(new_n1122), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1099), .A2(new_n1102), .B1(new_n1103), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1031), .B1(new_n984), .B2(new_n1032), .ZN(new_n1129));
  OAI21_X1  g704(.A(G286), .B1(new_n1036), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1039), .A2(new_n1033), .A3(G168), .A4(new_n1035), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(G8), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT51), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1131), .A2(new_n1134), .A3(G8), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1107), .A2(new_n1112), .A3(new_n1118), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1103), .B1(new_n1139), .B2(G301), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1133), .A2(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1055), .A2(new_n1128), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1015), .A2(new_n1016), .A3(new_n585), .A4(new_n589), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1009), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1013), .B(KEYINPUT113), .Z(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1050), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT62), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1135), .B1(new_n1132), .B2(KEYINPUT51), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1054), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1053), .A2(new_n1051), .A3(new_n1028), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n971), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT46), .B1(new_n958), .B2(new_n959), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT127), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(KEYINPUT127), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n963), .B(new_n785), .C1(new_n1166), .C2(G1996), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1164), .A2(new_n1165), .B1(new_n1167), .B2(new_n958), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT47), .Z(new_n1169));
  INV_X1    g744(.A(new_n958), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1170), .A2(G1986), .A3(G290), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT48), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n969), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n965), .A2(new_n967), .B1(new_n1071), .B2(new_n877), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT126), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1170), .B1(new_n1174), .B2(KEYINPUT126), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g753(.A1(new_n460), .A2(G227), .ZN(new_n1180));
  NOR3_X1   g754(.A1(G229), .A2(G401), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1181), .B1(new_n948), .B2(new_n942), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n902), .A2(new_n903), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1183), .ZN(G308));
  OAI221_X1 g758(.A(new_n1181), .B1(new_n902), .B2(new_n903), .C1(new_n942), .C2(new_n948), .ZN(G225));
endmodule


