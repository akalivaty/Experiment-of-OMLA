//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  INV_X1    g0022(.A(KEYINPUT69), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n222), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT67), .B(G238), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT68), .B(G77), .Z(new_n230));
  AOI22_X1  g0030(.A1(new_n229), .A2(G68), .B1(new_n230), .B2(G244), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n227), .B(new_n231), .C1(new_n223), .C2(new_n226), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n210), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n220), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT70), .ZN(new_n242));
  INV_X1    g0042(.A(G250), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT71), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n230), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(G1698), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT73), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n261), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G274), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n214), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n269), .ZN(new_n279));
  INV_X1    g0079(.A(new_n275), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n270), .A2(new_n275), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n276), .A2(new_n281), .B1(G226), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n272), .A2(G190), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT76), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n272), .A2(new_n284), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G200), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n208), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n208), .A2(new_n256), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT74), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(new_n294), .B1(G20), .B2(new_n204), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n294), .B2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n214), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n207), .A2(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G50), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n302), .A2(new_n305), .B1(new_n201), .B2(new_n301), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(KEYINPUT9), .A3(new_n306), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n288), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n286), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n285), .B(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n288), .A2(new_n309), .A3(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n287), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n272), .A2(new_n321), .A3(new_n284), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n307), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n230), .A2(G20), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n324), .B1(new_n292), .B2(new_n289), .C1(new_n290), .C2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n230), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n300), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n300), .A2(new_n328), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n326), .A2(new_n298), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n298), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G77), .A3(new_n303), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n276), .A2(new_n281), .ZN(new_n337));
  INV_X1    g0137(.A(G244), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n282), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n260), .A2(new_n239), .A3(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(G107), .B2(new_n260), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n266), .B2(new_n228), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n342), .B2(new_n271), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n336), .B1(new_n343), .B2(G190), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n343), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n343), .A2(new_n321), .B1(new_n335), .B2(new_n333), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n342), .A2(new_n271), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n319), .B1(new_n348), .B2(new_n339), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n318), .A2(new_n323), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n292), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(G58), .B(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G20), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT81), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n258), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G33), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(G20), .B1(new_n360), .B2(new_n257), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n257), .ZN(new_n364));
  AND2_X1   g0164(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g0165(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n367), .B2(G33), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n368), .A2(KEYINPUT7), .A3(G20), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n356), .C1(new_n363), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n362), .A2(G20), .ZN(new_n372));
  AOI21_X1  g0172(.A(G33), .B1(new_n358), .B2(new_n359), .ZN(new_n373));
  INV_X1    g0173(.A(new_n259), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n362), .B1(new_n262), .B2(G20), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n203), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n356), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n371), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n379), .A3(new_n298), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n274), .A2(new_n273), .A3(new_n275), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT72), .B1(new_n279), .B2(new_n280), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n381), .A2(new_n382), .B1(new_n239), .B2(new_n282), .ZN(new_n383));
  MUX2_X1   g0183(.A(G223), .B(G226), .S(G1698), .Z(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n360), .A3(new_n257), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n270), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n345), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n387), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n276), .A2(new_n281), .B1(G232), .B2(new_n283), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n289), .B1(new_n207), .B2(G20), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n302), .B1(new_n301), .B2(new_n289), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n380), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT17), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n380), .A2(new_n393), .A3(new_n398), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n380), .A2(new_n395), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n319), .B1(new_n383), .B2(new_n387), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n389), .A2(new_n390), .A3(new_n321), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT82), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n401), .A2(new_n405), .A3(new_n410), .A4(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n203), .A2(G20), .ZN(new_n413));
  INV_X1    g0213(.A(G77), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n290), .B2(new_n414), .C1(new_n201), .C2(new_n292), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n298), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n332), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT12), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n334), .B2(new_n303), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n420), .B1(KEYINPUT12), .B2(new_n301), .C1(new_n422), .C2(new_n203), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G226), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n239), .B2(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n262), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(KEYINPUT77), .A2(G33), .A3(G97), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n270), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(KEYINPUT78), .A3(new_n434), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n437), .A2(new_n438), .B1(G238), .B2(new_n283), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n337), .A2(KEYINPUT79), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n276), .A2(new_n442), .A3(new_n281), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n440), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n426), .B(G169), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(G179), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n450), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n426), .B1(new_n453), .B2(G169), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n425), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(G200), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n424), .C1(new_n391), .C2(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n352), .A2(new_n412), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n208), .A2(G87), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n368), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n260), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n208), .B2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n464), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(KEYINPUT24), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n464), .A2(new_n471), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n298), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n298), .B(new_n301), .C1(new_n207), .C2(G33), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT25), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n300), .B2(G107), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n300), .A2(new_n479), .A3(G107), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n478), .A2(G107), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT92), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n207), .B(G45), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(G264), .B(new_n270), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G257), .A2(G1698), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n243), .B2(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n360), .A2(new_n257), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G294), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n491), .B1(new_n496), .B2(new_n271), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n270), .A2(G274), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G1), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n488), .A2(G41), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(KEYINPUT84), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n485), .B1(new_n497), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n270), .B1(new_n494), .B2(new_n495), .ZN(new_n510));
  NOR4_X1   g0310(.A1(new_n510), .A2(new_n506), .A3(new_n491), .A4(KEYINPUT92), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(G169), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT93), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n497), .A2(new_n507), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n321), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n508), .A2(new_n511), .A3(new_n319), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT93), .B1(new_n519), .B2(new_n516), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n484), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n477), .A2(new_n483), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n391), .B1(new_n508), .B2(new_n511), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n515), .A2(new_n345), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G238), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n338), .B2(G1698), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n360), .A3(new_n257), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n270), .B1(new_n529), .B2(new_n465), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n503), .A2(new_n277), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n243), .B1(new_n502), .B2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n270), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n321), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n203), .A2(G20), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n360), .A2(new_n257), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n430), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n432), .A2(KEYINPUT19), .A3(new_n433), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n208), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n298), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n325), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n478), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n332), .A2(new_n325), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n319), .B1(new_n530), .B2(new_n534), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n536), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n478), .A2(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(new_n552), .A3(new_n548), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n530), .A2(G190), .A3(new_n534), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n345), .B1(new_n530), .B2(new_n534), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT88), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n545), .A2(new_n548), .ZN(new_n559));
  INV_X1    g0359(.A(new_n556), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n552), .C1(new_n560), .C2(new_n554), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n536), .A2(new_n549), .A3(new_n550), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT88), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n338), .A2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT4), .B1(new_n368), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G283), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n262), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  AND2_X1   g0373(.A1(G250), .A2(G1698), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(new_n262), .B2(new_n574), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n573), .A2(new_n257), .A3(new_n259), .A4(new_n574), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n271), .B1(new_n567), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G257), .B(new_n270), .C1(new_n487), .C2(new_n489), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n487), .A2(new_n500), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT84), .B1(new_n503), .B2(new_n504), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(new_n499), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n469), .B1(new_n375), .B2(new_n376), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  INV_X1    g0387(.A(G97), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n587), .A2(new_n588), .A3(G107), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n591), .A2(new_n208), .B1(new_n414), .B2(new_n292), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n298), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n300), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n478), .B2(G97), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n585), .A2(new_n319), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n578), .A2(new_n321), .A3(new_n584), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT86), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n360), .A2(new_n257), .A3(new_n566), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n257), .A2(new_n259), .A3(new_n574), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n262), .A2(new_n573), .A3(new_n574), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n606), .A3(new_n572), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n583), .B1(new_n607), .B2(new_n271), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n599), .B1(new_n608), .B2(new_n321), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n596), .B1(new_n598), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n593), .A2(new_n595), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n578), .A2(new_n391), .A3(new_n584), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n568), .B1(new_n260), .B2(new_n570), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n270), .B1(new_n615), .B2(new_n602), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n345), .B1(new_n616), .B2(new_n583), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n613), .ZN(new_n619));
  INV_X1    g0419(.A(new_n298), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n292), .A2(new_n414), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n590), .A2(new_n587), .ZN(new_n622));
  INV_X1    g0422(.A(new_n589), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n624), .B2(G20), .ZN(new_n625));
  INV_X1    g0425(.A(new_n372), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n256), .B1(new_n365), .B2(new_n366), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n259), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT7), .B1(new_n260), .B2(new_n208), .ZN(new_n629));
  OAI21_X1  g0429(.A(G107), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n620), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n478), .A2(G97), .ZN(new_n632));
  INV_X1    g0432(.A(new_n594), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT85), .B1(new_n619), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n610), .B1(new_n618), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n565), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n608), .A2(G169), .B1(new_n631), .B2(new_n634), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n608), .A2(new_n599), .A3(new_n321), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n616), .A2(G190), .A3(new_n583), .ZN(new_n644));
  AOI21_X1  g0444(.A(G200), .B1(new_n578), .B2(new_n584), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n635), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n611), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n619), .A2(KEYINPUT85), .A3(new_n635), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(G270), .B(new_n270), .C1(new_n487), .C2(new_n489), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n506), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(G264), .A2(G1698), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n245), .B2(G1698), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n360), .A2(new_n257), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(KEYINPUT89), .B(G303), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n260), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n271), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n345), .B1(new_n652), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G116), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n207), .B2(G33), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n620), .B(new_n662), .C1(new_n330), .C2(new_n331), .ZN(new_n663));
  INV_X1    g0463(.A(new_n331), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n661), .A3(new_n329), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n297), .A2(new_n214), .B1(G20), .B2(new_n661), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n568), .B(new_n208), .C1(G33), .C2(new_n588), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT20), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n666), .A2(KEYINPUT20), .A3(new_n667), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n663), .B(new_n665), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT90), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n650), .B1(new_n582), .B2(new_n499), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n270), .B1(new_n655), .B2(new_n657), .ZN(new_n673));
  OAI21_X1  g0473(.A(G200), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n670), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G190), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n671), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT21), .ZN(new_n681));
  OAI21_X1  g0481(.A(G169), .B1(new_n672), .B2(new_n673), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n675), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n652), .A2(new_n659), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n670), .A3(KEYINPUT21), .A4(G169), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n678), .A2(G179), .A3(new_n670), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT91), .B1(new_n680), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n671), .A2(new_n677), .A3(new_n679), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n649), .A2(KEYINPUT87), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n459), .A2(new_n526), .A3(new_n639), .A4(new_n693), .ZN(G372));
  INV_X1    g0494(.A(new_n323), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n409), .A2(new_n411), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n350), .ZN(new_n698));
  OAI21_X1  g0498(.A(G169), .B1(new_n445), .B2(new_n446), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT14), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n451), .A3(new_n447), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n457), .A2(new_n698), .B1(new_n701), .B2(new_n425), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n400), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n457), .A2(new_n698), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n705), .A2(new_n703), .A3(new_n455), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n697), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n695), .B1(new_n707), .B2(new_n318), .ZN(new_n708));
  INV_X1    g0508(.A(new_n459), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n647), .A2(new_n648), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n522), .B1(new_n519), .B2(new_n516), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n689), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n523), .A2(new_n524), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n557), .B1(new_n484), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT26), .B1(new_n643), .B2(new_n561), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n558), .A2(new_n643), .A3(KEYINPUT26), .A4(new_n564), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n551), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n708), .B1(new_n709), .B2(new_n719), .ZN(G369));
  NAND3_X1  g0520(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(KEYINPUT27), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT95), .Z(new_n723));
  INV_X1    g0523(.A(G213), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n721), .B2(KEYINPUT27), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G343), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n711), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n689), .A2(new_n728), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n526), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n728), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n526), .B1(new_n484), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n521), .A2(new_n728), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n675), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n688), .B2(new_n692), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n687), .A2(new_n736), .ZN(new_n738));
  OR3_X1    g0538(.A1(new_n737), .A2(KEYINPUT96), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT96), .B1(new_n737), .B2(new_n738), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n735), .A2(new_n739), .A3(G330), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n731), .B1(new_n743), .B2(new_n744), .ZN(G399));
  INV_X1    g0545(.A(new_n211), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G41), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n542), .A2(new_n661), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(G1), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n217), .B2(new_n748), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT29), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n719), .B2(new_n728), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT99), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT99), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n757), .B(new_n754), .C1(new_n719), .C2(new_n728), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n649), .B(new_n714), .C1(new_n521), .C2(new_n687), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n596), .B(new_n561), .C1(new_n598), .C2(new_n609), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n551), .B1(new_n760), .B2(KEYINPUT26), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT26), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n558), .A2(new_n643), .A3(new_n762), .A4(new_n564), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n728), .B1(new_n759), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT29), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n756), .A2(new_n758), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G330), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n693), .A2(new_n639), .A3(new_n526), .A4(new_n732), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n684), .A2(new_n321), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n535), .A2(new_n497), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n771), .A3(new_n608), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT98), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n678), .A2(new_n535), .A3(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n515), .A3(new_n585), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n770), .A2(new_n771), .A3(new_n608), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n728), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT31), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n768), .B1(new_n769), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n767), .A2(KEYINPUT100), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT100), .B1(new_n767), .B2(new_n784), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n753), .B1(new_n789), .B2(G1), .ZN(G364));
  AND2_X1   g0590(.A1(new_n208), .A2(G13), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G45), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n748), .A2(G1), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n739), .A2(new_n740), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n208), .A2(new_n321), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n803), .A2(new_n391), .A3(G200), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT103), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G58), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n208), .A2(G179), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n808), .A2(new_n391), .A3(G200), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT104), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G107), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n391), .A2(new_n345), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n808), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G87), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n802), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G190), .A2(G200), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n802), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G50), .A2(new_n817), .B1(new_n820), .B2(new_n230), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n807), .A2(new_n811), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n803), .A2(new_n345), .A3(G190), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n260), .B1(new_n823), .B2(G68), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n808), .A2(new_n818), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT32), .B1(new_n825), .B2(new_n353), .ZN(new_n826));
  OR3_X1    g0626(.A1(new_n825), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n391), .A2(G179), .A3(G200), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n208), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G97), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G326), .A2(new_n817), .B1(new_n820), .B2(G311), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n262), .B1(new_n814), .B2(G303), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n829), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT33), .B(G317), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n823), .A2(new_n837), .B1(new_n804), .B2(G322), .ZN(new_n838));
  INV_X1    g0638(.A(new_n825), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G329), .ZN(new_n840));
  INV_X1    g0640(.A(new_n810), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n822), .A2(new_n832), .B1(new_n836), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n214), .B1(G20), .B2(new_n319), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n799), .A2(new_n845), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT102), .Z(new_n848));
  NAND2_X1  g0648(.A1(new_n211), .A2(new_n262), .ZN(new_n849));
  INV_X1    g0649(.A(G355), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n850), .B1(G116), .B2(new_n211), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT101), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n746), .A2(new_n368), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(G45), .B2(new_n217), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n251), .B2(G45), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n848), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n846), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n794), .B1(new_n801), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n796), .A2(G330), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n795), .A2(new_n768), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n793), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT105), .Z(G396));
  NAND2_X1  g0663(.A1(new_n336), .A2(new_n728), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n346), .A2(new_n864), .B1(new_n347), .B2(new_n349), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n350), .A2(new_n728), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n719), .B2(new_n728), .ZN(new_n870));
  INV_X1    g0670(.A(new_n718), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n715), .B2(new_n716), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n351), .B(new_n732), .C1(new_n872), .C2(new_n551), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n794), .B1(new_n874), .B2(new_n784), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n784), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n845), .A2(new_n797), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n793), .B1(new_n414), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n869), .ZN(new_n879));
  INV_X1    g0679(.A(new_n845), .ZN(new_n880));
  INV_X1    g0680(.A(new_n823), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n881), .A2(new_n842), .B1(new_n469), .B2(new_n813), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G116), .B2(new_n820), .ZN(new_n883));
  INV_X1    g0683(.A(G303), .ZN(new_n884));
  INV_X1    g0684(.A(G311), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n816), .A2(new_n884), .B1(new_n825), .B2(new_n885), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n262), .B(new_n886), .C1(G294), .C2(new_n804), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n810), .A2(G87), .ZN(new_n888));
  AND4_X1   g0688(.A1(new_n831), .A2(new_n883), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n841), .A2(new_n203), .ZN(new_n890));
  AOI22_X1  g0690(.A1(G50), .A2(new_n814), .B1(new_n839), .B2(G132), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n368), .C1(new_n202), .C2(new_n829), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n823), .A2(G150), .B1(G159), .B2(new_n820), .ZN(new_n893));
  INV_X1    g0693(.A(G137), .ZN(new_n894));
  INV_X1    g0694(.A(G143), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n893), .B1(new_n894), .B2(new_n816), .C1(new_n805), .C2(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT34), .Z(new_n897));
  AOI211_X1 g0697(.A(new_n890), .B(new_n892), .C1(new_n897), .C2(KEYINPUT106), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n878), .B1(new_n879), .B2(new_n798), .C1(new_n880), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n876), .A2(new_n901), .ZN(G384));
  OR2_X1    g0702(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n216), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT36), .Z(new_n906));
  OAI211_X1 g0706(.A(new_n230), .B(new_n218), .C1(new_n202), .C2(new_n203), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n201), .A2(G68), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n207), .B(G13), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n873), .A2(new_n868), .ZN(new_n911));
  INV_X1    g0711(.A(new_n726), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n401), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n408), .A2(new_n913), .A3(new_n914), .A4(new_n396), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n370), .A2(new_n298), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT7), .B1(new_n368), .B2(G20), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n361), .A2(new_n362), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(G68), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT16), .B1(new_n919), .B2(new_n356), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n395), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n405), .A3(new_n407), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n912), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n922), .A2(new_n396), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n915), .B1(new_n924), .B2(new_n914), .ZN(new_n925));
  INV_X1    g0725(.A(new_n923), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n412), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n728), .B1(new_n419), .B2(new_n423), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT107), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n728), .C1(new_n419), .C2(new_n423), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n455), .A2(new_n457), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n701), .A2(new_n425), .A3(new_n728), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n911), .A2(new_n931), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n696), .A2(new_n726), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n701), .A2(new_n425), .A3(new_n732), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n400), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n397), .A2(KEYINPUT108), .A3(new_n399), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(new_n409), .A3(new_n411), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n913), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n408), .A2(new_n396), .A3(new_n913), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT37), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n948), .A2(new_n949), .B1(new_n915), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n944), .B(new_n930), .C1(new_n952), .C2(KEYINPUT38), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT38), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT39), .B1(new_n954), .B2(new_n928), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n943), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n942), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n756), .A2(new_n459), .A3(new_n758), .A4(new_n766), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n708), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n769), .A2(new_n782), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n869), .B1(new_n937), .B2(new_n938), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n954), .A2(new_n928), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n930), .B1(new_n952), .B2(KEYINPUT38), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n967), .A2(KEYINPUT40), .A3(new_n962), .A4(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n459), .A2(new_n962), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(G330), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n960), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n207), .B2(new_n791), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n960), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n910), .B1(new_n975), .B2(new_n976), .ZN(G367));
  OAI21_X1  g0777(.A(new_n847), .B1(new_n211), .B2(new_n325), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n246), .B2(new_n853), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n806), .A2(new_n656), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n881), .A2(new_n835), .B1(new_n825), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G283), .B2(new_n820), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n814), .A2(G116), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n984), .A2(new_n985), .B1(new_n469), .B2(new_n829), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n885), .A2(new_n816), .B1(new_n809), .B2(new_n588), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n368), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n980), .A2(new_n983), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n830), .A2(G68), .ZN(new_n991));
  INV_X1    g0791(.A(new_n804), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n291), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT110), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n823), .A2(G159), .B1(G50), .B2(new_n820), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT111), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n262), .B1(new_n825), .B2(new_n894), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n327), .A2(new_n809), .B1(new_n895), .B2(new_n816), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G58), .C2(new_n814), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n990), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n793), .B(new_n979), .C1(new_n1003), .C2(new_n845), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n728), .A2(new_n553), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n561), .A2(new_n562), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n551), .A2(new_n553), .A3(new_n728), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n799), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n792), .A2(G1), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n731), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n649), .B1(new_n635), .B2(new_n732), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n643), .A2(new_n728), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1016), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n731), .B2(new_n1014), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n731), .A2(new_n1014), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT45), .B1(new_n731), .B2(new_n1014), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1017), .B(new_n1019), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n743), .B2(new_n744), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT97), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n796), .A2(new_n1026), .A3(G330), .A4(new_n735), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1020), .B(new_n1021), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n742), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n526), .A2(new_n730), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n735), .B2(new_n730), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n860), .B(new_n1034), .Z(new_n1035));
  OAI22_X1  g0835(.A1(new_n1032), .A2(new_n1035), .B1(new_n786), .B2(new_n787), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n747), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1010), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1014), .A2(new_n526), .A3(new_n730), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT42), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n521), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n610), .B1(new_n1012), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1040), .A2(KEYINPUT42), .B1(new_n732), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1041), .A2(new_n1044), .B1(KEYINPUT43), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(KEYINPUT43), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1027), .A2(new_n742), .A3(new_n1014), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1009), .B1(new_n1039), .B2(new_n1050), .ZN(G387));
  NAND2_X1  g0851(.A1(new_n788), .A2(new_n1035), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1035), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n786), .B2(new_n787), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n747), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1010), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n240), .A2(G45), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n289), .A2(G50), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT50), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n750), .B(new_n502), .C1(new_n203), .C2(new_n414), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n853), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(G107), .B2(new_n211), .C1(new_n750), .C2(new_n849), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n793), .B1(new_n1062), .B2(new_n848), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n841), .A2(new_n588), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G159), .A2(new_n817), .B1(new_n820), .B2(G68), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n830), .A2(new_n546), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n368), .A3(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n881), .A2(new_n289), .B1(new_n825), .B2(new_n291), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n814), .A2(new_n230), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n992), .B2(new_n201), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G326), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n809), .A2(new_n661), .B1(new_n825), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n823), .A2(G311), .B1(new_n656), .B2(new_n820), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n816), .C1(new_n805), .C2(new_n981), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n830), .A2(G283), .B1(new_n814), .B2(G294), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n368), .B(new_n1073), .C1(new_n1082), .C2(KEYINPUT49), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(KEYINPUT49), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1071), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1063), .B1(new_n735), .B2(new_n800), .C1(new_n1085), .C2(new_n880), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1056), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1055), .A2(new_n1087), .ZN(G393));
  NAND3_X1  g0888(.A1(new_n1054), .A2(KEYINPUT115), .A3(new_n1032), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT115), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n767), .A2(new_n784), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT100), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1035), .B1(new_n1093), .B2(new_n785), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1090), .B1(new_n1094), .B2(new_n1031), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n747), .B1(new_n1054), .B2(new_n1032), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1015), .A2(new_n799), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT113), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n853), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n847), .B1(new_n588), .B2(new_n211), .C1(new_n1103), .C2(new_n254), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n794), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n804), .A2(G159), .B1(new_n817), .B2(G150), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI22_X1  g0907(.A1(new_n881), .A2(new_n201), .B1(new_n825), .B2(new_n895), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n203), .A2(new_n813), .B1(new_n819), .B2(new_n289), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n368), .B1(new_n414), .B2(new_n829), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n888), .A3(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n804), .A2(G311), .B1(new_n817), .B2(G317), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n823), .A2(new_n656), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n835), .B2(new_n819), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G283), .B2(new_n814), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n260), .B1(new_n825), .B2(new_n1075), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G116), .B2(new_n830), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1115), .A2(new_n811), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1113), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1105), .B1(new_n1123), .B2(new_n845), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1031), .A2(new_n1010), .B1(new_n1102), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1099), .A2(new_n1125), .ZN(G390));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n728), .B(new_n865), .C1(new_n759), .C2(new_n764), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n867), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n518), .A2(new_n520), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n687), .B1(new_n1130), .B2(new_n522), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n710), .A2(new_n610), .A3(new_n714), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n761), .A2(new_n763), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n732), .B(new_n866), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(KEYINPUT116), .A3(new_n868), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1129), .A2(new_n1136), .A3(new_n939), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n967), .A2(new_n943), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n939), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n873), .B2(new_n868), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n943), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n955), .B(new_n953), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n783), .A2(new_n963), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1140), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n953), .A2(new_n955), .A3(new_n797), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n793), .B1(new_n289), .B2(new_n877), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n881), .A2(new_n894), .B1(new_n819), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G159), .B2(new_n830), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT118), .Z(new_n1154));
  NOR2_X1   g0954(.A1(new_n813), .A2(new_n291), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n260), .B1(new_n839), .B2(G125), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n809), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(G50), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n804), .A2(G132), .B1(new_n817), .B2(G128), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G283), .A2(new_n817), .B1(new_n820), .B2(G97), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n469), .B2(new_n881), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT119), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n804), .A2(G116), .B1(G294), .B2(new_n839), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n260), .A3(new_n815), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1166), .B(new_n890), .C1(G77), .C2(new_n830), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1154), .A2(new_n1161), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1150), .B1(new_n1168), .B2(new_n880), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT120), .Z(new_n1170));
  AOI22_X1  g0970(.A1(new_n1148), .A2(new_n1010), .B1(new_n1149), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n459), .A2(new_n783), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n958), .A2(new_n708), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n962), .A2(G330), .A3(new_n879), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1141), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1176), .A3(new_n1145), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n939), .B1(new_n783), .B2(new_n879), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n962), .A2(new_n963), .A3(G330), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n911), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT117), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(new_n1148), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1127), .B(new_n867), .C1(new_n765), .C2(new_n866), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT116), .B1(new_n1135), .B2(new_n868), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1138), .B1(new_n1188), .B2(new_n939), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1143), .B1(new_n911), .B2(new_n939), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n953), .A2(new_n955), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1179), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1140), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT117), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n747), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1171), .B1(new_n1185), .B2(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(new_n877), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n794), .B1(G50), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n318), .A2(new_n323), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n307), .A2(new_n912), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT55), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n318), .A2(new_n323), .A3(new_n1203), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1208), .A3(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(new_n798), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n823), .B1(new_n804), .B2(G107), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n842), .B2(new_n825), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G116), .A2(new_n817), .B1(new_n820), .B2(new_n546), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n809), .A2(new_n202), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n991), .A3(new_n1069), .A4(new_n1218), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1215), .A2(new_n1219), .A3(G41), .A4(new_n368), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G50), .B1(new_n256), .B2(new_n486), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n368), .B2(G41), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n992), .A2(new_n1226), .B1(new_n813), .B2(new_n1151), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G125), .A2(new_n817), .B1(new_n820), .B2(G137), .ZN(new_n1228));
  INV_X1    g1028(.A(G132), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n881), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1227), .B(new_n1230), .C1(G150), .C2(new_n830), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT59), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT122), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1158), .A2(G159), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G33), .B(G41), .C1(new_n839), .C2(G124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(KEYINPUT122), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1225), .B1(KEYINPUT58), .B2(new_n1220), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1200), .B(new_n1213), .C1(new_n845), .C2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n966), .A2(G330), .A3(new_n968), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1212), .A2(new_n966), .A3(G330), .A4(new_n968), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n957), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n957), .A3(new_n1244), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1240), .B1(new_n1249), .B2(new_n1010), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n958), .A2(new_n708), .A3(new_n1172), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1148), .B2(new_n1181), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1243), .A2(new_n957), .A3(new_n1244), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n957), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n747), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1193), .A2(new_n1194), .A3(new_n1181), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1173), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1258), .B2(new_n1249), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1250), .B1(new_n1256), .B2(new_n1259), .ZN(G375));
  OAI22_X1  g1060(.A1(new_n881), .A2(new_n661), .B1(new_n819), .B2(new_n469), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G283), .B2(new_n804), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n816), .A2(new_n835), .B1(new_n813), .B2(new_n588), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n262), .B(new_n1263), .C1(G303), .C2(new_n839), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n810), .A2(G77), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1066), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n881), .A2(new_n1151), .B1(new_n819), .B2(new_n291), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1217), .B(new_n1267), .C1(G132), .C2(new_n817), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n806), .A2(G137), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n830), .A2(G50), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n368), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n813), .A2(new_n353), .B1(new_n825), .B2(new_n1226), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT124), .Z(new_n1273));
  OAI21_X1  g1073(.A(new_n1266), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n845), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1275), .B(new_n794), .C1(G68), .C2(new_n1199), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1141), .B2(new_n797), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1181), .B2(new_n1010), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1182), .A2(new_n1038), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(G381));
  OR2_X1    g1081(.A1(G381), .A2(G384), .ZN(new_n1282));
  INV_X1    g1082(.A(G396), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1055), .A3(new_n1087), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G390), .A2(new_n1282), .A3(G387), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1149), .A2(new_n1170), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1010), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1286), .B1(new_n1195), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n748), .B1(new_n1184), .B2(new_n1148), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(G375), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1285), .A2(new_n1291), .A3(new_n1292), .ZN(G407));
  NOR2_X1   g1093(.A1(new_n1285), .A2(new_n727), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1291), .ZN(new_n1295));
  OAI21_X1  g1095(.A(G213), .B1(new_n1294), .B2(new_n1295), .ZN(G409));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n724), .A2(G343), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1250), .C1(new_n1256), .C2(new_n1259), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1258), .A2(new_n1249), .A3(new_n1038), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1250), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1291), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1251), .A2(KEYINPUT60), .A3(new_n1180), .A4(new_n1177), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n747), .A4(new_n1182), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(G384), .A3(new_n1278), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1309), .B2(new_n1278), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1305), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1310), .A3(new_n1304), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1297), .B1(new_n1303), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(KEYINPUT126), .B(new_n1297), .C1(new_n1303), .C2(new_n1316), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1303), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT62), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1303), .A2(new_n1324), .A3(new_n1321), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1319), .A2(new_n1320), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G387), .A2(new_n1099), .A3(new_n1125), .ZN(new_n1327));
  XOR2_X1   g1127(.A(new_n1048), .B(new_n1049), .Z(new_n1328));
  AOI22_X1  g1128(.A1(new_n1053), .A2(new_n1031), .B1(new_n1093), .B2(new_n785), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1287), .B1(new_n1329), .B2(new_n1037), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1328), .A2(new_n1330), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1097), .B1(new_n1095), .B2(new_n1089), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1125), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1327), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT125), .B1(G390), .B2(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G393), .A2(G396), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1284), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1335), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1327), .A2(new_n1334), .A3(KEYINPUT125), .A4(new_n1338), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1326), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1317), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1322), .A2(KEYINPUT63), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1322), .A2(KEYINPUT63), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1345), .B(new_n1342), .C1(new_n1346), .C2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1344), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1291), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT125), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1334), .A2(new_n1351), .ZN(new_n1352));
  AOI22_X1  g1152(.A1(new_n1352), .A2(new_n1338), .B1(new_n1334), .B2(new_n1327), .ZN(new_n1353));
  AND4_X1   g1153(.A1(KEYINPUT125), .A2(new_n1327), .A3(new_n1334), .A4(new_n1338), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1299), .B(new_n1350), .C1(new_n1353), .C2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1350), .A2(new_n1299), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1340), .A2(new_n1341), .A3(new_n1356), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1355), .A2(new_n1321), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1321), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(G402));
endmodule


