

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n691, n692, n693,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727;

  INV_X1 U373 ( .A(n695), .ZN(n353) );
  INV_X1 U374 ( .A(n695), .ZN(n356) );
  AND2_X1 U375 ( .A1(n378), .A2(n415), .ZN(n604) );
  NAND2_X1 U376 ( .A1(n544), .A2(n352), .ZN(n380) );
  BUF_X1 U377 ( .A(n638), .Z(n351) );
  AND2_X1 U378 ( .A1(n372), .A2(n543), .ZN(n352) );
  XNOR2_X1 U379 ( .A(n369), .B(KEYINPUT39), .ZN(n554) );
  AND2_X1 U380 ( .A1(n571), .A2(n570), .ZN(n663) );
  XOR2_X1 U381 ( .A(KEYINPUT38), .B(n539), .Z(n623) );
  XNOR2_X1 U382 ( .A(n462), .B(n451), .ZN(n682) );
  XNOR2_X1 U383 ( .A(n709), .B(G146), .ZN(n462) );
  XNOR2_X1 U384 ( .A(G134), .B(G122), .ZN(n493) );
  XOR2_X1 U385 ( .A(G104), .B(G122), .Z(n502) );
  XOR2_X1 U386 ( .A(G116), .B(G107), .Z(n494) );
  XNOR2_X1 U387 ( .A(G119), .B(G110), .ZN(n466) );
  INV_X1 U388 ( .A(n604), .ZN(n711) );
  NAND2_X1 U389 ( .A1(n696), .A2(n604), .ZN(n652) );
  XNOR2_X2 U390 ( .A(n439), .B(n438), .ZN(n545) );
  NOR2_X2 U391 ( .A1(G953), .A2(n643), .ZN(n645) );
  AND2_X1 U392 ( .A1(n354), .A2(n353), .ZN(G63) );
  XNOR2_X1 U393 ( .A(n688), .B(n355), .ZN(n354) );
  INV_X1 U394 ( .A(n689), .ZN(n355) );
  AND2_X1 U395 ( .A1(n357), .A2(n356), .ZN(G66) );
  XNOR2_X1 U396 ( .A(n692), .B(n358), .ZN(n357) );
  INV_X1 U397 ( .A(n693), .ZN(n358) );
  INV_X2 U398 ( .A(KEYINPUT69), .ZN(n394) );
  XOR2_X1 U399 ( .A(G116), .B(G119), .Z(n454) );
  XNOR2_X1 U400 ( .A(G143), .B(G113), .ZN(n506) );
  XNOR2_X1 U401 ( .A(n576), .B(KEYINPUT33), .ZN(n639) );
  XNOR2_X2 U402 ( .A(n366), .B(KEYINPUT45), .ZN(n647) );
  XNOR2_X2 U403 ( .A(n394), .B(G131), .ZN(n503) );
  NOR2_X1 U404 ( .A1(n723), .A2(n725), .ZN(n536) );
  XOR2_X1 U405 ( .A(KEYINPUT4), .B(n491), .Z(n441) );
  XNOR2_X1 U406 ( .A(n409), .B(n371), .ZN(n592) );
  XNOR2_X1 U407 ( .A(n547), .B(n546), .ZN(n560) );
  XNOR2_X1 U408 ( .A(n442), .B(n441), .ZN(n709) );
  XNOR2_X1 U409 ( .A(n393), .B(n440), .ZN(n442) );
  XNOR2_X1 U410 ( .A(n503), .B(G137), .ZN(n393) );
  XNOR2_X1 U411 ( .A(n477), .B(n478), .ZN(n710) );
  XNOR2_X1 U412 ( .A(n428), .B(n429), .ZN(n457) );
  XNOR2_X1 U413 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U414 ( .A(n425), .B(KEYINPUT72), .ZN(n429) );
  INV_X2 U415 ( .A(G953), .ZN(n712) );
  XOR2_X1 U416 ( .A(KEYINPUT70), .B(G134), .Z(n440) );
  BUF_X2 U417 ( .A(n691), .Z(n359) );
  AND2_X2 U418 ( .A1(n421), .A2(n654), .ZN(n691) );
  NOR2_X2 U419 ( .A1(n583), .A2(n593), .ZN(n576) );
  NOR2_X2 U420 ( .A1(n560), .A2(n559), .ZN(n575) );
  NOR2_X1 U421 ( .A1(n570), .A2(n609), .ZN(n605) );
  INV_X1 U422 ( .A(G469), .ZN(n387) );
  NOR2_X1 U423 ( .A1(n674), .A2(n360), .ZN(n589) );
  OR2_X1 U424 ( .A1(G237), .A2(G902), .ZN(n516) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n379) );
  INV_X1 U426 ( .A(G472), .ZN(n405) );
  XNOR2_X1 U427 ( .A(n414), .B(KEYINPUT75), .ZN(n413) );
  INV_X1 U428 ( .A(KEYINPUT16), .ZN(n414) );
  XNOR2_X1 U429 ( .A(n383), .B(n382), .ZN(n687) );
  INV_X1 U430 ( .A(n710), .ZN(n382) );
  XNOR2_X1 U431 ( .A(n511), .B(n384), .ZN(n383) );
  XNOR2_X1 U432 ( .A(n510), .B(n508), .ZN(n384) );
  XNOR2_X1 U433 ( .A(G110), .B(KEYINPUT73), .ZN(n443) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(KEYINPUT94), .Z(n444) );
  XOR2_X1 U435 ( .A(G101), .B(G140), .Z(n445) );
  XOR2_X1 U436 ( .A(G104), .B(G107), .Z(n448) );
  NAND2_X1 U437 ( .A1(n541), .A2(n623), .ZN(n369) );
  AND2_X1 U438 ( .A1(n562), .A2(n368), .ZN(n563) );
  AND2_X1 U439 ( .A1(n593), .A2(n570), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n575), .B(KEYINPUT0), .ZN(n585) );
  AND2_X1 U441 ( .A1(n605), .A2(n406), .ZN(n588) );
  INV_X1 U442 ( .A(KEYINPUT22), .ZN(n371) );
  AND2_X1 U443 ( .A1(n561), .A2(n411), .ZN(n410) );
  NAND2_X1 U444 ( .A1(n691), .A2(G475), .ZN(n392) );
  NAND2_X1 U445 ( .A1(n691), .A2(G210), .ZN(n402) );
  NOR2_X1 U446 ( .A1(n667), .A2(n627), .ZN(n552) );
  INV_X1 U447 ( .A(n726), .ZN(n373) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n484) );
  XOR2_X1 U449 ( .A(G902), .B(KEYINPUT89), .Z(n437) );
  NOR2_X1 U450 ( .A1(G953), .A2(G237), .ZN(n458) );
  INV_X1 U451 ( .A(KEYINPUT3), .ZN(n426) );
  XOR2_X1 U452 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n507) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n432) );
  XNOR2_X1 U454 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n397), .B(KEYINPUT18), .ZN(n396) );
  NAND2_X1 U456 ( .A1(n712), .A2(G224), .ZN(n397) );
  INV_X1 U457 ( .A(n609), .ZN(n411) );
  XNOR2_X1 U458 ( .A(n575), .B(KEYINPUT0), .ZN(n412) );
  NOR2_X1 U459 ( .A1(n677), .A2(n416), .ZN(n415) );
  XNOR2_X1 U460 ( .A(n380), .B(n379), .ZN(n378) );
  INV_X1 U461 ( .A(n676), .ZN(n416) );
  XOR2_X1 U462 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n478) );
  INV_X1 U463 ( .A(KEYINPUT1), .ZN(n452) );
  NOR2_X1 U464 ( .A1(n668), .A2(n528), .ZN(n517) );
  AND2_X1 U465 ( .A1(n535), .A2(n534), .ZN(n541) );
  AND2_X1 U466 ( .A1(n588), .A2(n403), .ZN(n534) );
  BUF_X1 U467 ( .A(n545), .Z(n539) );
  INV_X1 U468 ( .A(KEYINPUT19), .ZN(n546) );
  XNOR2_X1 U469 ( .A(n529), .B(n367), .ZN(n530) );
  INV_X1 U470 ( .A(KEYINPUT28), .ZN(n367) );
  NOR2_X1 U471 ( .A1(n584), .A2(n528), .ZN(n529) );
  NAND2_X1 U472 ( .A1(n691), .A2(G472), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n466), .B(n413), .ZN(n424) );
  INV_X1 U474 ( .A(KEYINPUT121), .ZN(n374) );
  XNOR2_X1 U475 ( .A(n408), .B(n407), .ZN(n723) );
  INV_X1 U476 ( .A(KEYINPUT40), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n566), .B(n565), .ZN(n722) );
  XNOR2_X1 U478 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n565) );
  NOR2_X1 U479 ( .A1(n567), .A2(n564), .ZN(n566) );
  NAND2_X1 U480 ( .A1(n537), .A2(n381), .ZN(n668) );
  INV_X1 U481 ( .A(n550), .ZN(n381) );
  OR2_X1 U482 ( .A1(n548), .A2(n560), .ZN(n667) );
  NAND2_X1 U483 ( .A1(n588), .A2(n584), .ZN(n398) );
  INV_X1 U484 ( .A(KEYINPUT60), .ZN(n389) );
  INV_X1 U485 ( .A(KEYINPUT56), .ZN(n399) );
  NOR2_X1 U486 ( .A1(n587), .A2(n398), .ZN(n360) );
  XNOR2_X1 U487 ( .A(n483), .B(KEYINPUT25), .ZN(n594) );
  AND2_X1 U488 ( .A1(n642), .A2(n641), .ZN(n361) );
  XOR2_X1 U489 ( .A(n656), .B(KEYINPUT62), .Z(n362) );
  XNOR2_X1 U490 ( .A(KEYINPUT66), .B(n651), .ZN(n363) );
  XOR2_X1 U491 ( .A(n687), .B(n686), .Z(n364) );
  XNOR2_X1 U492 ( .A(n680), .B(n679), .ZN(n365) );
  INV_X1 U493 ( .A(n695), .ZN(n418) );
  NAND2_X1 U494 ( .A1(n652), .A2(KEYINPUT82), .ZN(n377) );
  NAND2_X1 U495 ( .A1(n602), .A2(n603), .ZN(n366) );
  XNOR2_X1 U496 ( .A(n375), .B(n374), .ZN(n643) );
  NOR2_X1 U497 ( .A1(n373), .A2(n553), .ZN(n372) );
  XNOR2_X1 U498 ( .A(n648), .B(KEYINPUT83), .ZN(n386) );
  OR2_X2 U499 ( .A1(n652), .A2(n653), .ZN(n421) );
  NOR2_X1 U500 ( .A1(n594), .A2(n609), .ZN(n490) );
  NAND2_X1 U501 ( .A1(n370), .A2(n590), .ZN(n597) );
  XNOR2_X1 U502 ( .A(n589), .B(KEYINPUT99), .ZN(n370) );
  NAND2_X1 U503 ( .A1(n385), .A2(n363), .ZN(n654) );
  INV_X1 U504 ( .A(n592), .ZN(n567) );
  NAND2_X1 U505 ( .A1(n592), .A2(n568), .ZN(n569) );
  XNOR2_X1 U506 ( .A(n392), .B(n364), .ZN(n391) );
  NAND2_X1 U507 ( .A1(n391), .A2(n418), .ZN(n390) );
  NAND2_X1 U508 ( .A1(n581), .A2(n582), .ZN(n599) );
  XNOR2_X1 U509 ( .A(n390), .B(n389), .ZN(G60) );
  NAND2_X1 U510 ( .A1(n386), .A2(n604), .ZN(n385) );
  NAND2_X1 U511 ( .A1(n376), .A2(n361), .ZN(n375) );
  XNOR2_X1 U512 ( .A(n377), .B(KEYINPUT2), .ZN(n376) );
  INV_X1 U513 ( .A(n537), .ZN(n549) );
  INV_X1 U514 ( .A(n668), .ZN(n670) );
  XNOR2_X2 U515 ( .A(n533), .B(n452), .ZN(n606) );
  XNOR2_X2 U516 ( .A(n388), .B(n387), .ZN(n533) );
  OR2_X2 U517 ( .A1(n682), .A2(G902), .ZN(n388) );
  XNOR2_X2 U518 ( .A(KEYINPUT71), .B(G101), .ZN(n427) );
  NAND2_X1 U519 ( .A1(n412), .A2(n410), .ZN(n409) );
  NOR2_X1 U520 ( .A1(n655), .A2(G902), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n400), .B(n399), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n401), .A2(n418), .ZN(n400) );
  XNOR2_X1 U523 ( .A(n402), .B(n365), .ZN(n401) );
  XNOR2_X1 U524 ( .A(n404), .B(n532), .ZN(n403) );
  NAND2_X1 U525 ( .A1(n615), .A2(n622), .ZN(n404) );
  XNOR2_X2 U526 ( .A(n463), .B(n405), .ZN(n615) );
  INV_X1 U527 ( .A(n533), .ZN(n406) );
  NAND2_X1 U528 ( .A1(n554), .A2(n670), .ZN(n408) );
  XNOR2_X1 U529 ( .A(n417), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U530 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U531 ( .A(n420), .B(n362), .ZN(n419) );
  XNOR2_X1 U532 ( .A(n569), .B(KEYINPUT65), .ZN(n571) );
  NOR2_X1 U533 ( .A1(G952), .A2(n712), .ZN(n695) );
  XNOR2_X1 U534 ( .A(n462), .B(n461), .ZN(n655) );
  XNOR2_X1 U535 ( .A(n441), .B(n432), .ZN(n435) );
  NOR2_X1 U536 ( .A1(n582), .A2(n572), .ZN(n574) );
  XNOR2_X1 U537 ( .A(n457), .B(n456), .ZN(n460) );
  XNOR2_X1 U538 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U540 ( .A(KEYINPUT87), .ZN(n524) );
  XNOR2_X1 U541 ( .A(n585), .B(KEYINPUT93), .ZN(n587) );
  XNOR2_X1 U542 ( .A(n424), .B(n423), .ZN(n431) );
  BUF_X1 U543 ( .A(n647), .Z(n696) );
  XNOR2_X1 U544 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n606), .B(n524), .ZN(n562) );
  XNOR2_X1 U546 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U547 ( .A(n594), .ZN(n570) );
  XNOR2_X1 U548 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U549 ( .A(n494), .B(n502), .Z(n423) );
  XNOR2_X2 U550 ( .A(G113), .B(KEYINPUT90), .ZN(n425) );
  XNOR2_X1 U551 ( .A(n457), .B(KEYINPUT74), .ZN(n430) );
  XNOR2_X1 U552 ( .A(n430), .B(n431), .ZN(n705) );
  XOR2_X2 U553 ( .A(G143), .B(G128), .Z(n491) );
  XOR2_X1 U554 ( .A(G146), .B(G125), .Z(n476) );
  XNOR2_X1 U555 ( .A(KEYINPUT73), .B(n476), .ZN(n433) );
  XOR2_X1 U556 ( .A(n433), .B(KEYINPUT86), .Z(n434) );
  XNOR2_X1 U557 ( .A(n705), .B(n436), .ZN(n678) );
  XNOR2_X1 U558 ( .A(KEYINPUT15), .B(n437), .ZN(n646) );
  NAND2_X1 U559 ( .A1(n678), .A2(n646), .ZN(n439) );
  AND2_X1 U560 ( .A1(G210), .A2(n516), .ZN(n438) );
  XNOR2_X1 U561 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U562 ( .A(n446), .B(n445), .ZN(n450) );
  NAND2_X1 U563 ( .A1(G227), .A2(n712), .ZN(n447) );
  XNOR2_X1 U564 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U565 ( .A(KEYINPUT5), .B(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U566 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U567 ( .A(n455), .B(KEYINPUT97), .Z(n456) );
  XOR2_X1 U568 ( .A(KEYINPUT77), .B(n458), .Z(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(G210), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n615), .B(KEYINPUT6), .ZN(n593) );
  NAND2_X1 U571 ( .A1(G234), .A2(n646), .ZN(n464) );
  XNOR2_X1 U572 ( .A(KEYINPUT20), .B(n464), .ZN(n480) );
  NAND2_X1 U573 ( .A1(G221), .A2(n480), .ZN(n465) );
  XNOR2_X1 U574 ( .A(KEYINPUT21), .B(n465), .ZN(n609) );
  XNOR2_X1 U575 ( .A(G128), .B(G137), .ZN(n467) );
  XNOR2_X1 U576 ( .A(n467), .B(n466), .ZN(n471) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n469) );
  XNOR2_X1 U578 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n468) );
  XNOR2_X1 U579 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U580 ( .A(n471), .B(n470), .ZN(n475) );
  NAND2_X1 U581 ( .A1(n712), .A2(G234), .ZN(n473) );
  XNOR2_X1 U582 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n473), .B(n472), .ZN(n492) );
  NAND2_X1 U584 ( .A1(n492), .A2(G221), .ZN(n474) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n476), .B(G140), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n479), .B(n710), .ZN(n693) );
  NOR2_X1 U588 ( .A1(G902), .A2(n693), .ZN(n482) );
  NAND2_X1 U589 ( .A1(G217), .A2(n480), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n484), .B(KEYINPUT14), .ZN(n485) );
  XNOR2_X1 U592 ( .A(KEYINPUT76), .B(n485), .ZN(n487) );
  NAND2_X1 U593 ( .A1(G902), .A2(n487), .ZN(n556) );
  NOR2_X1 U594 ( .A1(G900), .A2(n556), .ZN(n486) );
  NAND2_X1 U595 ( .A1(G953), .A2(n486), .ZN(n489) );
  NAND2_X1 U596 ( .A1(n487), .A2(G952), .ZN(n488) );
  XNOR2_X1 U597 ( .A(n488), .B(KEYINPUT91), .ZN(n635) );
  NAND2_X1 U598 ( .A1(n635), .A2(n712), .ZN(n555) );
  NAND2_X1 U599 ( .A1(n489), .A2(n555), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n490), .A2(n535), .ZN(n528) );
  XNOR2_X1 U601 ( .A(n491), .B(KEYINPUT104), .ZN(n500) );
  NAND2_X1 U602 ( .A1(n492), .A2(G217), .ZN(n498) );
  XNOR2_X1 U603 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U605 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U606 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n500), .B(n499), .ZN(n689) );
  NOR2_X1 U608 ( .A1(G902), .A2(n689), .ZN(n501) );
  XOR2_X1 U609 ( .A(G478), .B(n501), .Z(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n505) );
  XNOR2_X1 U611 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n505), .B(n504), .ZN(n511) );
  XNOR2_X1 U613 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U614 ( .A1(G214), .A2(n509), .ZN(n510) );
  NOR2_X1 U615 ( .A1(n687), .A2(G902), .ZN(n515) );
  XOR2_X1 U616 ( .A(KEYINPUT13), .B(KEYINPUT102), .Z(n513) );
  XNOR2_X1 U617 ( .A(KEYINPUT103), .B(G475), .ZN(n512) );
  XNOR2_X1 U618 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U619 ( .A(n515), .B(n514), .ZN(n537) );
  NAND2_X1 U620 ( .A1(G214), .A2(n516), .ZN(n622) );
  NAND2_X1 U621 ( .A1(n517), .A2(n622), .ZN(n518) );
  NOR2_X1 U622 ( .A1(n593), .A2(n518), .ZN(n522) );
  XNOR2_X1 U623 ( .A(KEYINPUT107), .B(n522), .ZN(n519) );
  NOR2_X1 U624 ( .A1(n606), .A2(n519), .ZN(n520) );
  XNOR2_X1 U625 ( .A(n520), .B(KEYINPUT43), .ZN(n521) );
  NOR2_X1 U626 ( .A1(n539), .A2(n521), .ZN(n677) );
  AND2_X1 U627 ( .A1(n539), .A2(n522), .ZN(n523) );
  XNOR2_X1 U628 ( .A(KEYINPUT36), .B(n523), .ZN(n525) );
  NAND2_X1 U629 ( .A1(n525), .A2(n562), .ZN(n526) );
  XNOR2_X1 U630 ( .A(n526), .B(KEYINPUT110), .ZN(n726) );
  NAND2_X1 U631 ( .A1(n623), .A2(n622), .ZN(n628) );
  NOR2_X1 U632 ( .A1(n537), .A2(n550), .ZN(n561) );
  INV_X1 U633 ( .A(n561), .ZN(n625) );
  NOR2_X1 U634 ( .A1(n628), .A2(n625), .ZN(n527) );
  XNOR2_X1 U635 ( .A(KEYINPUT41), .B(n527), .ZN(n638) );
  INV_X1 U636 ( .A(n615), .ZN(n584) );
  OR2_X1 U637 ( .A1(n530), .A2(n533), .ZN(n548) );
  NOR2_X1 U638 ( .A1(n638), .A2(n548), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n531), .B(KEYINPUT42), .ZN(n725) );
  XOR2_X1 U640 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n532) );
  XNOR2_X1 U641 ( .A(n536), .B(KEYINPUT46), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n537), .A2(n550), .ZN(n538) );
  XOR2_X1 U643 ( .A(n538), .B(KEYINPUT106), .Z(n578) );
  AND2_X1 U644 ( .A1(n539), .A2(n578), .ZN(n540) );
  NAND2_X1 U645 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U646 ( .A(KEYINPUT109), .B(n542), .ZN(n720) );
  INV_X1 U647 ( .A(n720), .ZN(n543) );
  NAND2_X1 U648 ( .A1(n545), .A2(n622), .ZN(n547) );
  NAND2_X1 U649 ( .A1(n550), .A2(n549), .ZN(n664) );
  NAND2_X1 U650 ( .A1(n664), .A2(n668), .ZN(n551) );
  XNOR2_X1 U651 ( .A(KEYINPUT105), .B(n551), .ZN(n627) );
  XOR2_X1 U652 ( .A(KEYINPUT47), .B(n552), .Z(n553) );
  INV_X1 U653 ( .A(n664), .ZN(n673) );
  NAND2_X1 U654 ( .A1(n554), .A2(n673), .ZN(n676) );
  INV_X1 U655 ( .A(n555), .ZN(n558) );
  XOR2_X1 U656 ( .A(KEYINPUT92), .B(G898), .Z(n700) );
  NAND2_X1 U657 ( .A1(G953), .A2(n700), .ZN(n704) );
  NOR2_X1 U658 ( .A1(n556), .A2(n704), .ZN(n557) );
  NOR2_X1 U659 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U660 ( .A(n563), .B(KEYINPUT81), .ZN(n564) );
  INV_X1 U661 ( .A(n606), .ZN(n591) );
  AND2_X1 U662 ( .A1(n584), .A2(n591), .ZN(n568) );
  NOR2_X1 U663 ( .A1(n722), .A2(n663), .ZN(n582) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n572) );
  INV_X1 U665 ( .A(KEYINPUT64), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n574), .B(n573), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n605), .A2(n606), .ZN(n583) );
  NOR2_X1 U668 ( .A1(n587), .A2(n639), .ZN(n577) );
  XNOR2_X1 U669 ( .A(n577), .B(KEYINPUT34), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X2 U671 ( .A(n580), .B(KEYINPUT35), .ZN(n721) );
  NOR2_X1 U672 ( .A1(n721), .A2(KEYINPUT44), .ZN(n581) );
  NOR2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n618) );
  NAND2_X1 U674 ( .A1(n585), .A2(n618), .ZN(n586) );
  XNOR2_X1 U675 ( .A(n586), .B(KEYINPUT31), .ZN(n674) );
  INV_X1 U676 ( .A(n627), .ZN(n590) );
  AND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n596) );
  AND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n657) );
  AND2_X1 U680 ( .A1(n597), .A2(n657), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n601) );
  AND2_X1 U682 ( .A1(n721), .A2(KEYINPUT44), .ZN(n600) );
  NOR2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U684 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n608) );
  OR2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n608), .B(n607), .ZN(n613) );
  XOR2_X1 U687 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n611) );
  NAND2_X1 U688 ( .A1(n609), .A2(n570), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT116), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT51), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT117), .B(n620), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n351), .A2(n621), .ZN(n633) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n626), .B(KEYINPUT118), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U702 ( .A1(n631), .A2(n639), .ZN(n632) );
  NOR2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U704 ( .A(KEYINPUT52), .B(n634), .Z(n636) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U706 ( .A(KEYINPUT119), .B(n637), .Z(n642) );
  NOR2_X1 U707 ( .A1(n639), .A2(n351), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT120), .B(n640), .Z(n641) );
  XNOR2_X1 U709 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n645), .B(n644), .ZN(G75) );
  INV_X1 U711 ( .A(n646), .ZN(n649) );
  NAND2_X1 U712 ( .A1(n647), .A2(n649), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n649), .B(KEYINPUT84), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n653) );
  XOR2_X1 U716 ( .A(n655), .B(KEYINPUT111), .Z(n656) );
  XNOR2_X1 U717 ( .A(G101), .B(n657), .ZN(G3) );
  NAND2_X1 U718 ( .A1(n670), .A2(n360), .ZN(n658) );
  XNOR2_X1 U719 ( .A(G104), .B(n658), .ZN(G6) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .ZN(n662) );
  XOR2_X1 U721 ( .A(KEYINPUT26), .B(KEYINPUT112), .Z(n660) );
  NAND2_X1 U722 ( .A1(n360), .A2(n673), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U724 ( .A(n662), .B(n661), .ZN(G9) );
  XOR2_X1 U725 ( .A(n663), .B(G110), .Z(G12) );
  NOR2_X1 U726 ( .A1(n664), .A2(n667), .ZN(n666) );
  XNOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .ZN(n665) );
  XNOR2_X1 U728 ( .A(n666), .B(n665), .ZN(G30) );
  NOR2_X1 U729 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U730 ( .A(G146), .B(n669), .Z(G48) );
  XOR2_X1 U731 ( .A(G113), .B(KEYINPUT113), .Z(n672) );
  NAND2_X1 U732 ( .A1(n674), .A2(n670), .ZN(n671) );
  XNOR2_X1 U733 ( .A(n672), .B(n671), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n675), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(G134), .B(n676), .ZN(G36) );
  XOR2_X1 U737 ( .A(G140), .B(n677), .Z(G42) );
  XNOR2_X1 U738 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT85), .ZN(n679) );
  NAND2_X1 U740 ( .A1(n359), .A2(G469), .ZN(n684) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  NOR2_X1 U742 ( .A1(n695), .A2(n685), .ZN(G54) );
  XOR2_X1 U743 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n686) );
  NAND2_X1 U744 ( .A1(G478), .A2(n359), .ZN(n688) );
  NAND2_X1 U745 ( .A1(G217), .A2(n359), .ZN(n692) );
  NAND2_X1 U746 ( .A1(n696), .A2(n712), .ZN(n703) );
  NAND2_X1 U747 ( .A1(G224), .A2(G953), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n697), .B(KEYINPUT61), .ZN(n698) );
  XNOR2_X1 U749 ( .A(n698), .B(KEYINPUT123), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U751 ( .A(KEYINPUT124), .B(n701), .Z(n702) );
  NAND2_X1 U752 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U753 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U754 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U755 ( .A(KEYINPUT125), .B(n708), .ZN(G69) );
  XNOR2_X1 U756 ( .A(n709), .B(n710), .ZN(n714) );
  XNOR2_X1 U757 ( .A(n711), .B(n714), .ZN(n713) );
  NAND2_X1 U758 ( .A1(n713), .A2(n712), .ZN(n718) );
  XNOR2_X1 U759 ( .A(G227), .B(n714), .ZN(n715) );
  NAND2_X1 U760 ( .A1(n715), .A2(G900), .ZN(n716) );
  NAND2_X1 U761 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U762 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U763 ( .A(KEYINPUT126), .B(n719), .ZN(G72) );
  XOR2_X1 U764 ( .A(G143), .B(n720), .Z(G45) );
  XOR2_X1 U765 ( .A(n721), .B(G122), .Z(G24) );
  XOR2_X1 U766 ( .A(n722), .B(G119), .Z(G21) );
  XNOR2_X1 U767 ( .A(G131), .B(KEYINPUT127), .ZN(n724) );
  XNOR2_X1 U768 ( .A(n724), .B(n723), .ZN(G33) );
  XOR2_X1 U769 ( .A(n725), .B(G137), .Z(G39) );
  XOR2_X1 U770 ( .A(G125), .B(n726), .Z(n727) );
  XNOR2_X1 U771 ( .A(KEYINPUT37), .B(n727), .ZN(G27) );
endmodule

