

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n400), .B(n399), .ZN(n550) );
  XOR2_X1 U324 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n445) );
  XOR2_X1 U325 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n292) );
  XNOR2_X1 U326 ( .A(G71GAT), .B(G57GAT), .ZN(n291) );
  XNOR2_X1 U327 ( .A(n292), .B(n291), .ZN(n347) );
  XOR2_X1 U328 ( .A(KEYINPUT73), .B(G78GAT), .Z(n294) );
  XNOR2_X1 U329 ( .A(G148GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U330 ( .A(n294), .B(n293), .ZN(n421) );
  XNOR2_X1 U331 ( .A(n347), .B(n421), .ZN(n306) );
  XOR2_X1 U332 ( .A(G99GAT), .B(G85GAT), .Z(n337) );
  XOR2_X1 U333 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n296) );
  XNOR2_X1 U334 ( .A(G120GAT), .B(KEYINPUT75), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U336 ( .A(n337), .B(n297), .Z(n299) );
  NAND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U339 ( .A(n300), .B(KEYINPUT32), .ZN(n304) );
  XOR2_X1 U340 ( .A(G204GAT), .B(G64GAT), .Z(n302) );
  XNOR2_X1 U341 ( .A(G176GAT), .B(G92GAT), .ZN(n301) );
  XNOR2_X1 U342 ( .A(n302), .B(n301), .ZN(n401) );
  XOR2_X1 U343 ( .A(n401), .B(KEYINPUT31), .Z(n303) );
  XNOR2_X1 U344 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U345 ( .A(n306), .B(n305), .ZN(n573) );
  XOR2_X1 U346 ( .A(G22GAT), .B(G8GAT), .Z(n308) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G197GAT), .ZN(n307) );
  XNOR2_X1 U348 ( .A(n308), .B(n307), .ZN(n327) );
  XOR2_X1 U349 ( .A(G15GAT), .B(G1GAT), .Z(n354) );
  XOR2_X1 U350 ( .A(n354), .B(G36GAT), .Z(n316) );
  INV_X1 U351 ( .A(G43GAT), .ZN(n309) );
  NAND2_X1 U352 ( .A1(G29GAT), .A2(n309), .ZN(n312) );
  INV_X1 U353 ( .A(G29GAT), .ZN(n310) );
  NAND2_X1 U354 ( .A1(n310), .A2(G43GAT), .ZN(n311) );
  NAND2_X1 U355 ( .A1(n312), .A2(n311), .ZN(n314) );
  XNOR2_X1 U356 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n314), .B(n313), .ZN(n332) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(n332), .ZN(n315) );
  XNOR2_X1 U359 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U360 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n318) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U362 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U363 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U364 ( .A(KEYINPUT29), .B(G113GAT), .Z(n322) );
  XNOR2_X1 U365 ( .A(KEYINPUT69), .B(G141GAT), .ZN(n321) );
  XNOR2_X1 U366 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U367 ( .A(n323), .B(KEYINPUT30), .ZN(n324) );
  XNOR2_X1 U368 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U369 ( .A(n327), .B(n326), .ZN(n504) );
  NAND2_X1 U370 ( .A1(n573), .A2(n504), .ZN(n459) );
  XOR2_X1 U371 ( .A(KEYINPUT76), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U372 ( .A(KEYINPUT11), .B(KEYINPUT77), .ZN(n328) );
  XNOR2_X1 U373 ( .A(n329), .B(n328), .ZN(n344) );
  XOR2_X1 U374 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n331) );
  XNOR2_X1 U375 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n330) );
  XNOR2_X1 U376 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U377 ( .A(n332), .B(KEYINPUT65), .ZN(n334) );
  AND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U379 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U380 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U381 ( .A(G106GAT), .B(G218GAT), .Z(n339) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G190GAT), .Z(n410) );
  XNOR2_X1 U383 ( .A(n410), .B(n337), .ZN(n338) );
  XNOR2_X1 U384 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U385 ( .A(G50GAT), .B(G162GAT), .Z(n417) );
  XOR2_X1 U386 ( .A(n340), .B(n417), .Z(n341) );
  XNOR2_X1 U387 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U388 ( .A(n344), .B(n343), .Z(n538) );
  INV_X1 U389 ( .A(n538), .ZN(n561) );
  XOR2_X1 U390 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n346) );
  XNOR2_X1 U391 ( .A(G64GAT), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U392 ( .A(n346), .B(n345), .ZN(n358) );
  XOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .Z(n409) );
  XOR2_X1 U394 ( .A(n347), .B(n409), .Z(n349) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U396 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U397 ( .A(G78GAT), .B(KEYINPUT15), .Z(n351) );
  XNOR2_X1 U398 ( .A(G127GAT), .B(KEYINPUT78), .ZN(n350) );
  XNOR2_X1 U399 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U400 ( .A(n353), .B(n352), .Z(n356) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XNOR2_X1 U402 ( .A(n354), .B(n425), .ZN(n355) );
  XNOR2_X1 U403 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U404 ( .A(n358), .B(n357), .ZN(n578) );
  NOR2_X1 U405 ( .A1(n561), .A2(n578), .ZN(n359) );
  XOR2_X1 U406 ( .A(KEYINPUT79), .B(n359), .Z(n360) );
  XNOR2_X1 U407 ( .A(KEYINPUT16), .B(n360), .ZN(n443) );
  XOR2_X1 U408 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n362) );
  XNOR2_X1 U409 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n361) );
  XNOR2_X1 U410 ( .A(n362), .B(n361), .ZN(n379) );
  XOR2_X1 U411 ( .A(G155GAT), .B(G85GAT), .Z(n364) );
  XNOR2_X1 U412 ( .A(G29GAT), .B(G162GAT), .ZN(n363) );
  XNOR2_X1 U413 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U414 ( .A(KEYINPUT5), .B(G148GAT), .Z(n366) );
  XNOR2_X1 U415 ( .A(G1GAT), .B(G57GAT), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U417 ( .A(n368), .B(n367), .Z(n377) );
  XOR2_X1 U418 ( .A(G127GAT), .B(G134GAT), .Z(n370) );
  XNOR2_X1 U419 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n369) );
  XNOR2_X1 U420 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U421 ( .A(G113GAT), .B(n371), .Z(n394) );
  XNOR2_X1 U422 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n372), .B(KEYINPUT2), .ZN(n416) );
  XOR2_X1 U424 ( .A(n416), .B(KEYINPUT1), .Z(n374) );
  NAND2_X1 U425 ( .A1(G225GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n394), .B(n375), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U429 ( .A(n379), .B(n378), .Z(n546) );
  XOR2_X1 U430 ( .A(G183GAT), .B(G176GAT), .Z(n381) );
  XNOR2_X1 U431 ( .A(G15GAT), .B(G99GAT), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U433 ( .A(G43GAT), .B(G190GAT), .Z(n382) );
  XNOR2_X1 U434 ( .A(n383), .B(n382), .ZN(n398) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n385) );
  XNOR2_X1 U436 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U438 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n387) );
  XNOR2_X1 U439 ( .A(KEYINPUT82), .B(KEYINPUT64), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U441 ( .A(n389), .B(n388), .Z(n396) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n390), .B(KEYINPUT84), .ZN(n391) );
  XOR2_X1 U444 ( .A(n391), .B(KEYINPUT19), .Z(n393) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n413) );
  XNOR2_X1 U447 ( .A(n413), .B(n394), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n398), .B(n397), .ZN(n400) );
  NAND2_X1 U450 ( .A1(G227GAT), .A2(G233GAT), .ZN(n399) );
  XOR2_X1 U451 ( .A(KEYINPUT91), .B(n401), .Z(n403) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U453 ( .A(n403), .B(n402), .ZN(n408) );
  XNOR2_X1 U454 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n404), .B(KEYINPUT87), .ZN(n405) );
  XOR2_X1 U456 ( .A(n405), .B(KEYINPUT88), .Z(n407) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(G218GAT), .ZN(n406) );
  XNOR2_X1 U458 ( .A(n407), .B(n406), .ZN(n429) );
  XOR2_X1 U459 ( .A(n408), .B(n429), .Z(n412) );
  XNOR2_X1 U460 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U461 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U462 ( .A(n414), .B(n413), .ZN(n541) );
  XNOR2_X1 U463 ( .A(n541), .B(KEYINPUT27), .ZN(n415) );
  XNOR2_X1 U464 ( .A(KEYINPUT92), .B(n415), .ZN(n438) );
  XNOR2_X1 U465 ( .A(KEYINPUT68), .B(KEYINPUT28), .ZN(n430) );
  XOR2_X1 U466 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U467 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U468 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U469 ( .A(n420), .B(KEYINPUT23), .Z(n423) );
  XNOR2_X1 U470 ( .A(n421), .B(KEYINPUT22), .ZN(n422) );
  XNOR2_X1 U471 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U472 ( .A(n424), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U473 ( .A(n425), .B(G204GAT), .ZN(n426) );
  XNOR2_X1 U474 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U475 ( .A(n429), .B(n428), .ZN(n547) );
  XOR2_X1 U476 ( .A(n430), .B(n547), .Z(n489) );
  INV_X1 U477 ( .A(n489), .ZN(n431) );
  NAND2_X1 U478 ( .A1(n438), .A2(n431), .ZN(n509) );
  NOR2_X1 U479 ( .A1(n550), .A2(n509), .ZN(n432) );
  NOR2_X1 U480 ( .A1(n546), .A2(n432), .ZN(n442) );
  INV_X1 U481 ( .A(n546), .ZN(n526) );
  NAND2_X1 U482 ( .A1(n550), .A2(n541), .ZN(n433) );
  NAND2_X1 U483 ( .A1(n547), .A2(n433), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT25), .B(n434), .Z(n439) );
  NOR2_X1 U485 ( .A1(n550), .A2(n547), .ZN(n436) );
  XNOR2_X1 U486 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U488 ( .A(KEYINPUT93), .B(n437), .Z(n567) );
  NAND2_X1 U489 ( .A1(n567), .A2(n438), .ZN(n525) );
  NAND2_X1 U490 ( .A1(n439), .A2(n525), .ZN(n440) );
  NOR2_X1 U491 ( .A1(n526), .A2(n440), .ZN(n441) );
  NOR2_X1 U492 ( .A1(n442), .A2(n441), .ZN(n455) );
  NAND2_X1 U493 ( .A1(n443), .A2(n455), .ZN(n471) );
  NOR2_X1 U494 ( .A1(n459), .A2(n471), .ZN(n450) );
  NAND2_X1 U495 ( .A1(n450), .A2(n526), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(n446), .ZN(G1324GAT) );
  NAND2_X1 U498 ( .A1(n541), .A2(n450), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n447), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U500 ( .A(G15GAT), .B(KEYINPUT35), .Z(n449) );
  NAND2_X1 U501 ( .A1(n450), .A2(n550), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(G1326GAT) );
  NAND2_X1 U503 ( .A1(n450), .A2(n489), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U505 ( .A(KEYINPUT96), .B(KEYINPUT99), .Z(n453) );
  XNOR2_X1 U506 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n462) );
  XNOR2_X1 U508 ( .A(KEYINPUT36), .B(KEYINPUT97), .ZN(n454) );
  XOR2_X1 U509 ( .A(n454), .B(n538), .Z(n581) );
  NAND2_X1 U510 ( .A1(n455), .A2(n578), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n581), .A2(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT37), .B(KEYINPUT98), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n458), .B(n457), .ZN(n483) );
  NOR2_X1 U514 ( .A1(n459), .A2(n483), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT38), .ZN(n468) );
  NAND2_X1 U516 ( .A1(n468), .A2(n526), .ZN(n461) );
  XOR2_X1 U517 ( .A(n462), .B(n461), .Z(G1328GAT) );
  NAND2_X1 U518 ( .A1(n468), .A2(n541), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U520 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n467) );
  XOR2_X1 U521 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n465) );
  NAND2_X1 U522 ( .A1(n550), .A2(n468), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(G1330GAT) );
  XNOR2_X1 U525 ( .A(G50GAT), .B(KEYINPUT102), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n489), .A2(n468), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(G1331GAT) );
  XNOR2_X1 U528 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n473) );
  INV_X1 U529 ( .A(n504), .ZN(n569) );
  XNOR2_X1 U530 ( .A(n573), .B(KEYINPUT41), .ZN(n515) );
  NAND2_X1 U531 ( .A1(n569), .A2(n515), .ZN(n482) );
  NOR2_X1 U532 ( .A1(n482), .A2(n471), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n478), .A2(n526), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(G1332GAT) );
  XOR2_X1 U535 ( .A(G64GAT), .B(KEYINPUT103), .Z(n475) );
  NAND2_X1 U536 ( .A1(n478), .A2(n541), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n475), .B(n474), .ZN(G1333GAT) );
  NAND2_X1 U538 ( .A1(n478), .A2(n550), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT104), .ZN(n477) );
  XNOR2_X1 U540 ( .A(G71GAT), .B(n477), .ZN(G1334GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n480) );
  NAND2_X1 U542 ( .A1(n478), .A2(n489), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U544 ( .A(G78GAT), .B(n481), .Z(G1335GAT) );
  XNOR2_X1 U545 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n483), .A2(n482), .ZN(n490) );
  NAND2_X1 U547 ( .A1(n490), .A2(n526), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(G1336GAT) );
  XOR2_X1 U549 ( .A(G92GAT), .B(KEYINPUT107), .Z(n487) );
  NAND2_X1 U550 ( .A1(n490), .A2(n541), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(G1337GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n550), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n488), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n492) );
  NAND2_X1 U555 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U557 ( .A(G106GAT), .B(n493), .Z(G1339GAT) );
  AND2_X1 U558 ( .A1(n526), .A2(n550), .ZN(n511) );
  NAND2_X1 U559 ( .A1(n504), .A2(n515), .ZN(n494) );
  XNOR2_X1 U560 ( .A(KEYINPUT46), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(KEYINPUT109), .B(n578), .ZN(n558) );
  NOR2_X1 U562 ( .A1(n561), .A2(n558), .ZN(n495) );
  NAND2_X1 U563 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U564 ( .A(KEYINPUT47), .B(n497), .ZN(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT110), .B(n498), .ZN(n507) );
  NOR2_X1 U566 ( .A1(n578), .A2(n581), .ZN(n501) );
  XOR2_X1 U567 ( .A(KEYINPUT111), .B(KEYINPUT45), .Z(n499) );
  XNOR2_X1 U568 ( .A(KEYINPUT66), .B(n499), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(n502) );
  NAND2_X1 U570 ( .A1(n573), .A2(n502), .ZN(n503) );
  NOR2_X1 U571 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(KEYINPUT112), .B(n505), .ZN(n506) );
  NOR2_X1 U573 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT48), .B(n508), .ZN(n543) );
  NOR2_X1 U575 ( .A1(n543), .A2(n509), .ZN(n510) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n569), .A2(n518), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G113GAT), .B(n514), .ZN(G1340GAT) );
  INV_X1 U581 ( .A(n515), .ZN(n553) );
  NOR2_X1 U582 ( .A1(n553), .A2(n518), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n520) );
  INV_X1 U586 ( .A(n518), .ZN(n522) );
  NAND2_X1 U587 ( .A1(n522), .A2(n558), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(n521), .ZN(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n561), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  NOR2_X1 U593 ( .A1(n543), .A2(n525), .ZN(n527) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n569), .A2(n537), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G141GAT), .B(n529), .ZN(G1344GAT) );
  NOR2_X1 U598 ( .A1(n537), .A2(n553), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n531) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  NOR2_X1 U603 ( .A1(n578), .A2(n537), .ZN(n535) );
  XNOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  NOR2_X1 U607 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U608 ( .A(G162GAT), .B(n539), .Z(n540) );
  XNOR2_X1 U609 ( .A(KEYINPUT120), .B(n540), .ZN(G1347GAT) );
  XNOR2_X1 U610 ( .A(KEYINPUT121), .B(n541), .ZN(n542) );
  NOR2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(KEYINPUT54), .B(n544), .ZN(n545) );
  AND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n568) );
  NAND2_X1 U614 ( .A1(n568), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT122), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT55), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n569), .A2(n557), .ZN(n552) );
  XOR2_X1 U619 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n557), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n556), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n560) );
  INV_X1 U625 ( .A(n557), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n569), .A2(n580), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n580), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

