//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252;
  XOR2_X1   g0000(.A(KEYINPUT65), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND3_X1  g0004(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n218), .B(new_n219), .C1(new_n204), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n208), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n203), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n212), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(new_n233));
  NOR2_X1   g0033(.A1(new_n207), .A2(new_n223), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n217), .B(new_n230), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n227), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  INV_X1    g0041(.A(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n223), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n203), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT77), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT17), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT16), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n204), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G58), .A2(G68), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n205), .A2(new_n206), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G159), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n256), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT74), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT73), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n262), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n261), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n257), .A3(new_n212), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n262), .A2(G33), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n276), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT7), .B1(new_n283), .B2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G68), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n272), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT16), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n231), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT74), .B(new_n256), .C1(new_n266), .C2(new_n272), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n275), .A2(new_n287), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(new_n212), .A3(G1), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n289), .B1(new_n211), .B2(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT76), .ZN(new_n300));
  OR2_X1    g0100(.A1(G223), .A2(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n224), .A2(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n279), .A2(new_n261), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n260), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n211), .B(G274), .C1(G41), .C2(G45), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n312), .A2(new_n313), .B1(new_n315), .B2(new_n227), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n309), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT75), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n307), .B1(new_n303), .B2(new_n304), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n316), .ZN(new_n321));
  AOI21_X1  g0121(.A(G200), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n320), .A2(G190), .A3(new_n316), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n300), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT75), .B1(new_n309), .B2(new_n317), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n320), .A2(new_n319), .A3(new_n316), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n323), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(KEYINPUT76), .A3(new_n329), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n255), .B(new_n299), .C1(new_n324), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n330), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n291), .A2(new_n298), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT17), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n254), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT76), .B1(new_n328), .B2(new_n329), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n322), .A2(new_n300), .A3(new_n323), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n255), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n299), .B1(new_n324), .B2(new_n330), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(KEYINPUT77), .A3(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n320), .A2(G179), .A3(new_n316), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n318), .A2(new_n321), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n299), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n299), .A2(KEYINPUT18), .A3(new_n346), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n295), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n212), .A2(G33), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n289), .B1(new_n208), .B2(new_n293), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n297), .A2(G77), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n315), .A2(new_n225), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n312), .A2(new_n313), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G107), .ZN(new_n364));
  INV_X1    g0164(.A(G1698), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n258), .A2(new_n365), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n363), .B1(new_n364), .B2(new_n258), .C1(new_n366), .C2(new_n227), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n361), .B(new_n362), .C1(new_n367), .C2(new_n308), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n360), .B1(G190), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n325), .B2(new_n368), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n335), .A2(new_n342), .A3(new_n351), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n227), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G226), .B2(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G97), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n264), .B1(new_n260), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n362), .B1(new_n375), .B2(new_n308), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n220), .B2(new_n315), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n384), .A3(G169), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n270), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n387), .A2(new_n223), .B1(new_n212), .B2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n354), .A2(new_n208), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n289), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT11), .ZN(new_n391));
  OR3_X1    g0191(.A1(new_n294), .A2(KEYINPUT12), .A3(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT12), .B1(new_n294), .B2(G68), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(G68), .B2(new_n297), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n368), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n360), .C1(G169), .C2(new_n368), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n380), .A2(G200), .ZN(new_n400));
  INV_X1    g0200(.A(new_n395), .ZN(new_n401));
  INV_X1    g0201(.A(G190), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n380), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n294), .A2(new_n223), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n297), .B2(new_n223), .ZN(new_n406));
  XOR2_X1   g0206(.A(new_n406), .B(KEYINPUT71), .Z(new_n407));
  AOI21_X1  g0207(.A(new_n212), .B1(new_n201), .B2(new_n207), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n295), .A2(new_n354), .B1(new_n409), .B2(new_n387), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n289), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT9), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(G222), .ZN(new_n418));
  OR3_X1    g0218(.A1(new_n366), .A2(KEYINPUT69), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n264), .A2(G77), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT69), .B1(new_n366), .B2(new_n418), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n308), .ZN(new_n424));
  INV_X1    g0224(.A(new_n362), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n307), .A2(G226), .A3(new_n314), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G200), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n402), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n416), .A2(new_n417), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT10), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n427), .A2(G179), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n427), .A2(new_n345), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n436));
  AND4_X1   g0236(.A1(new_n414), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n371), .A2(new_n404), .A3(new_n432), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT86), .ZN(new_n439));
  OR2_X1    g0239(.A1(G257), .A2(G1698), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n365), .A2(G264), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n279), .A2(new_n261), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n264), .A2(G303), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n439), .B1(new_n444), .B2(new_n308), .ZN(new_n445));
  AOI211_X1 g0245(.A(KEYINPUT86), .B(new_n307), .C1(new_n442), .C2(new_n443), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G274), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n307), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n242), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n345), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n212), .C1(G33), .C2(new_n374), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT80), .B(G116), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n289), .B(new_n460), .C1(new_n461), .C2(new_n212), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT20), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n289), .B(new_n293), .C1(new_n211), .C2(G33), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(G116), .ZN(new_n467));
  INV_X1    g0267(.A(new_n461), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n293), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n458), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n444), .A2(new_n308), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n444), .A2(new_n439), .A3(new_n308), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n457), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G200), .ZN(new_n478));
  INV_X1    g0278(.A(new_n470), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n479), .C1(new_n402), .C2(new_n477), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(KEYINPUT21), .A3(G169), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n447), .A2(G179), .A3(new_n457), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT87), .B1(new_n483), .B2(new_n470), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT87), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n485), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n473), .B(new_n480), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n277), .B1(new_n262), .B2(G33), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n260), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n261), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n261), .A2(new_n263), .A3(G250), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n365), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n492), .A2(new_n495), .A3(new_n459), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n308), .ZN(new_n498));
  INV_X1    g0298(.A(new_n455), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G257), .B1(G274), .B2(new_n453), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n345), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n466), .A2(G97), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n294), .A2(G97), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n509), .A3(G107), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n510), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n507), .A2(new_n509), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(KEYINPUT79), .C1(new_n512), .C2(new_n511), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n212), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n387), .A2(new_n208), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n364), .B1(new_n259), .B2(new_n265), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n289), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n503), .B(new_n505), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n498), .A2(new_n500), .A3(new_n397), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n502), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n501), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n402), .C2(new_n501), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n487), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n279), .A2(G250), .A3(new_n365), .A4(new_n261), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT89), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT89), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n283), .A2(new_n535), .A3(G250), .A4(new_n365), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n537), .A2(KEYINPUT90), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n308), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n499), .A2(G264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n454), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(G190), .A3(new_n454), .A4(new_n545), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n466), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n293), .A2(new_n364), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT25), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n279), .A2(KEYINPUT22), .A3(G87), .A4(new_n261), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n461), .A2(G33), .ZN(new_n553));
  AOI21_X1  g0353(.A(G20), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n258), .A2(new_n212), .A3(G87), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT88), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT23), .ZN(new_n561));
  OAI211_X1 g0361(.A(G20), .B(new_n364), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT24), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NOR4_X1   g0367(.A1(new_n554), .A2(new_n558), .A3(new_n564), .A4(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n551), .B1(new_n569), .B2(new_n289), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n546), .A2(new_n345), .ZN(new_n572));
  OR3_X1    g0372(.A1(new_n566), .A2(new_n523), .A3(new_n568), .ZN(new_n573));
  INV_X1    g0373(.A(new_n551), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n549), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n544), .A2(new_n397), .A3(new_n454), .A4(new_n545), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n204), .A2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n279), .A2(new_n261), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT83), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n354), .B2(new_n374), .ZN(new_n582));
  NAND3_X1  g0382(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n212), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n374), .A3(new_n364), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(KEYINPUT82), .A3(new_n212), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n283), .A2(new_n591), .A3(new_n578), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n580), .A2(new_n582), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n590), .A2(new_n582), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT84), .A3(new_n580), .A4(new_n592), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n289), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n466), .A2(new_n355), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n356), .A2(new_n293), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G238), .A2(G1698), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n225), .B2(G1698), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n283), .A2(new_n603), .B1(G33), .B2(new_n461), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n449), .A2(G250), .ZN(new_n605));
  INV_X1    g0405(.A(G274), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n449), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n307), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n604), .A2(new_n307), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n345), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  INV_X1    g0411(.A(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n397), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(KEYINPUT81), .A3(new_n397), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n601), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n598), .A2(new_n600), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n609), .A2(G200), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n466), .A2(G87), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n609), .A2(new_n402), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n598), .A2(new_n600), .A3(new_n619), .A4(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT85), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n577), .A2(new_n616), .A3(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n438), .A2(new_n532), .A3(new_n571), .A4(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n396), .A2(new_n399), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n403), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n335), .A2(new_n342), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n351), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT92), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n432), .B(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n437), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n613), .A2(new_n610), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n601), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n526), .A4(new_n616), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n526), .B(new_n637), .C1(new_n622), .C2(new_n624), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT91), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n638), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n616), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n624), .B(new_n618), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n623), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n526), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n470), .A2(new_n483), .B1(new_n471), .B2(new_n472), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n577), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n531), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n637), .B1(new_n622), .B2(new_n624), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n571), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n643), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n438), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n635), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n648), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n292), .A2(G20), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n231), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT93), .ZN(new_n661));
  INV_X1    g0461(.A(G213), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n659), .B2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(KEYINPUT93), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n479), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n487), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n577), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n575), .A2(new_n667), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n571), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n577), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NOR4_X1   g0478(.A1(new_n445), .A2(new_n446), .A3(new_n397), .A4(new_n456), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n458), .B2(KEYINPUT21), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n485), .B1(new_n680), .B2(new_n479), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n483), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n667), .B1(new_n683), .B2(new_n473), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n674), .B1(new_n677), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n215), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n588), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n234), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n683), .A2(new_n577), .A3(new_n473), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n548), .A2(new_n570), .A3(new_n549), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n651), .B1(new_n697), .B2(new_n547), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n698), .A3(new_n650), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n646), .A2(new_n641), .A3(new_n526), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n699), .A2(new_n637), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n695), .B1(new_n702), .B2(new_n668), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n654), .A2(new_n695), .A3(new_n668), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n532), .A2(new_n627), .A3(new_n571), .A4(new_n668), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n544), .A2(new_n545), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n501), .A2(new_n609), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n679), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n679), .A4(new_n707), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n498), .B2(new_n500), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n546), .A2(new_n477), .A3(new_n609), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n667), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI211_X1 g0518(.A(new_n703), .B(new_n704), .C1(new_n718), .C2(G330), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n694), .B1(new_n719), .B2(G1), .ZN(G364));
  XNOR2_X1  g0520(.A(new_n672), .B(KEYINPUT94), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n658), .A2(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n689), .A2(G1), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT95), .Z(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n722), .B(new_n726), .C1(G330), .C2(new_n671), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n231), .B1(G20), .B2(new_n345), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n212), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G159), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT32), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n212), .A2(new_n402), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n397), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(new_n740), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n203), .B1(new_n742), .B2(new_n208), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT96), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n325), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n587), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n738), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n212), .A2(new_n397), .A3(new_n325), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n402), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n750), .A2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n748), .B1(new_n223), .B2(new_n752), .C1(new_n204), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n730), .A2(G190), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n374), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n745), .A2(new_n731), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n364), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n755), .A2(new_n264), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  INV_X1    g0563(.A(new_n741), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n753), .A2(new_n763), .B1(new_n764), .B2(G322), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT100), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n751), .A2(G326), .ZN(new_n767));
  INV_X1    g0567(.A(new_n742), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G311), .ZN(new_n769));
  INV_X1    g0569(.A(G303), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n264), .B1(new_n746), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  INV_X1    g0574(.A(G294), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n735), .A2(new_n774), .B1(new_n775), .B2(new_n758), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n760), .A2(new_n778), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n728), .B1(new_n762), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n687), .A2(new_n264), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G355), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n248), .A2(new_n448), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n687), .A2(new_n283), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n692), .B2(G45), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(G116), .B2(new_n215), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n728), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n726), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n781), .B(new_n792), .C1(new_n671), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n727), .A2(new_n794), .ZN(G396));
  OAI21_X1  g0595(.A(new_n283), .B1(new_n204), .B2(new_n760), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n753), .A2(G150), .B1(new_n751), .B2(G137), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT101), .Z(new_n798));
  INV_X1    g0598(.A(G143), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n799), .B2(new_n741), .C1(new_n736), .C2(new_n742), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT34), .Z(new_n801));
  INV_X1    g0601(.A(new_n746), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n796), .B(new_n801), .C1(G50), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n203), .B2(new_n758), .C1(new_n804), .C2(new_n735), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n264), .B1(new_n754), .B2(new_n778), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n760), .A2(new_n587), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n461), .B2(new_n768), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n770), .B2(new_n752), .C1(new_n758), .C2(new_n374), .ZN(new_n809));
  INV_X1    g0609(.A(new_n735), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n806), .B(new_n809), .C1(G311), .C2(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n364), .B2(new_n746), .C1(new_n775), .C2(new_n741), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n726), .B1(new_n813), .B2(new_n728), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n728), .A2(new_n788), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n360), .A2(new_n667), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n370), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n399), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n399), .A2(new_n667), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n814), .B1(G77), .B2(new_n816), .C1(new_n789), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n718), .A2(G330), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n654), .A2(new_n668), .A3(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n821), .B1(new_n654), .B2(new_n668), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n823), .B(new_n827), .Z(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n828), .B2(new_n725), .ZN(G384));
  NAND3_X1  g0629(.A1(new_n339), .A2(new_n351), .A3(new_n341), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n333), .A2(new_n665), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT104), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n347), .B1(new_n333), .B2(new_n665), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n340), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT37), .B1(new_n831), .B2(KEYINPUT103), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n833), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n335), .A2(new_n342), .A3(new_n351), .ZN(new_n843));
  INV_X1    g0643(.A(new_n665), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n287), .A2(new_n289), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT16), .B1(new_n285), .B2(new_n286), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n298), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n346), .B2(new_n844), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n338), .A2(new_n849), .ZN(new_n850));
  MUX2_X1   g0650(.A(new_n837), .B(new_n850), .S(KEYINPUT37), .Z(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n386), .A2(new_n395), .A3(new_n668), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n848), .A2(new_n851), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n841), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n852), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n852), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n403), .B1(new_n401), .B2(new_n668), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n396), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n856), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n824), .B2(new_n820), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n349), .A2(new_n350), .A3(new_n665), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n438), .B1(new_n704), .B2(new_n703), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n635), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n438), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n864), .A2(new_n821), .A3(new_n856), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n716), .A2(new_n717), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n853), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT40), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n862), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n873), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n853), .B2(new_n875), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n716), .A2(new_n878), .A3(new_n874), .A4(new_n717), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n852), .B2(new_n859), .ZN(new_n883));
  OAI21_X1  g0683(.A(G330), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n438), .A2(G330), .A3(new_n716), .A4(new_n717), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n880), .A2(new_n718), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n872), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n211), .B2(new_n658), .ZN(new_n888));
  INV_X1    g0688(.A(G116), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n516), .A2(new_n518), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(KEYINPUT35), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n233), .C1(KEYINPUT35), .C2(new_n890), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n234), .A2(G77), .A3(new_n267), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT102), .Z(new_n895));
  INV_X1    g0695(.A(new_n201), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n204), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G1), .A3(new_n292), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n893), .A3(new_n898), .ZN(G367));
  OAI21_X1  g0699(.A(new_n650), .B1(new_n528), .B2(new_n668), .ZN(new_n900));
  AND4_X1   g0700(.A1(new_n524), .A2(new_n502), .A3(new_n525), .A4(new_n667), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n677), .A3(new_n684), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT42), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n674), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n908), .B(new_n909), .C1(new_n527), .C2(new_n667), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n668), .B1(new_n617), .B2(new_n620), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n638), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n651), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT106), .Z(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n678), .A2(new_n905), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT107), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(KEYINPUT107), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n917), .B1(new_n916), .B2(new_n919), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n688), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n685), .A2(new_n906), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT45), .Z(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n685), .A2(new_n906), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(KEYINPUT44), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT44), .B2(new_n932), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n932), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n678), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT109), .B1(new_n677), .B2(new_n684), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n677), .A2(new_n684), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n939), .B(new_n940), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n672), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n722), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n719), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n928), .B1(new_n945), .B2(new_n719), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n723), .A2(G1), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n925), .B(new_n926), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n746), .A2(new_n949), .A3(new_n889), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n802), .A2(new_n461), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n283), .B1(new_n951), .B2(new_n949), .ZN(new_n952));
  INV_X1    g0752(.A(G311), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n752), .A2(new_n953), .B1(new_n770), .B2(new_n741), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n952), .B1(new_n775), .B2(new_n754), .C1(new_n954), .C2(KEYINPUT111), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n950), .B(new_n955), .C1(KEYINPUT111), .C2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(new_n760), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(G97), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n757), .A2(G107), .B1(G283), .B2(new_n768), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT110), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G317), .B2(new_n810), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n758), .A2(new_n204), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n760), .A2(new_n208), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n810), .B2(G137), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n752), .A2(new_n799), .B1(new_n201), .B2(new_n742), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G58), .B2(new_n802), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(new_n409), .C2(new_n741), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n963), .B(new_n968), .C1(G159), .C2(new_n753), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n962), .B1(new_n258), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n728), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n913), .A2(new_n793), .ZN(new_n974));
  INV_X1    g0774(.A(new_n785), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n791), .B1(new_n215), .B2(new_n356), .C1(new_n243), .C2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n725), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n948), .A2(new_n977), .ZN(G387));
  AND2_X1   g0778(.A1(new_n943), .A2(new_n947), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT113), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n689), .B1(new_n943), .B2(new_n719), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n719), .B2(new_n943), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n280), .B1(new_n468), .B2(new_n760), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G317), .A2(new_n764), .B1(new_n768), .B2(G303), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT114), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n953), .B2(new_n754), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G322), .B2(new_n751), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT48), .Z(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n778), .B2(new_n758), .C1(new_n775), .C2(new_n746), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT49), .Z(new_n990));
  AOI211_X1 g0790(.A(new_n983), .B(new_n990), .C1(G326), .C2(new_n810), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n758), .A2(new_n356), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G159), .B2(new_n751), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n958), .C1(new_n409), .C2(new_n735), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n280), .B(new_n994), .C1(G50), .C2(new_n764), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n802), .A2(G77), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n753), .A2(new_n352), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G68), .B2(new_n768), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n728), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n975), .B1(new_n239), .B2(G45), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n690), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n782), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n352), .A2(new_n223), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n204), .A2(new_n208), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1005), .A2(G45), .A3(new_n1006), .A4(new_n1002), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1003), .A2(new_n1007), .B1(G107), .B2(new_n215), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n726), .B1(new_n1008), .B2(new_n791), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1000), .B(new_n1009), .C1(new_n677), .C2(new_n793), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n980), .A2(new_n982), .A3(new_n1010), .ZN(G393));
  AOI21_X1  g0811(.A(new_n689), .B1(new_n938), .B2(new_n944), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n945), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n791), .B1(new_n975), .B2(new_n252), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G97), .B2(new_n687), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n757), .A2(G77), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n751), .A2(G150), .B1(G159), .B2(new_n764), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(KEYINPUT51), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n283), .B1(new_n746), .B2(new_n204), .C1(new_n754), .C2(new_n201), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n807), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n799), .B2(new_n735), .C1(new_n295), .C2(new_n742), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n264), .B1(new_n746), .B2(new_n778), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n751), .A2(G317), .B1(G311), .B2(new_n764), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n761), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n770), .B2(new_n754), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(G322), .C2(new_n810), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(KEYINPUT52), .B2(new_n1024), .C1(new_n775), .C2(new_n742), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n758), .A2(new_n468), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1022), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n726), .B(new_n1015), .C1(new_n1030), .C2(new_n728), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n906), .B2(new_n793), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n947), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n938), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1013), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G390));
  NAND2_X1  g0836(.A1(new_n855), .A2(new_n860), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n824), .A2(new_n820), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n865), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT115), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n856), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT115), .B1(new_n866), .B2(new_n857), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n702), .A2(new_n668), .A3(new_n819), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1045), .A2(new_n820), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n853), .B(new_n856), .C1(new_n1046), .C2(new_n865), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n716), .A2(G330), .A3(new_n717), .A4(new_n821), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n865), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n718), .A2(G330), .A3(new_n821), .A4(new_n1039), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1044), .A2(new_n1052), .A3(new_n1047), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n947), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1037), .A2(new_n788), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n810), .A2(G125), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n757), .A2(G159), .B1(G128), .B2(new_n751), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n258), .B1(new_n201), .B2(new_n760), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT54), .B(G143), .Z(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n742), .B1(new_n804), .B2(new_n741), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1058), .B(new_n1061), .C1(G137), .C2(new_n753), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n746), .A2(new_n409), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT53), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1056), .A2(new_n1057), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n264), .B1(new_n752), .B2(new_n778), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n747), .B(new_n1066), .C1(G116), .C2(new_n764), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n810), .A2(G294), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n753), .A2(G107), .B1(G68), .B2(new_n957), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1067), .A2(new_n1016), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n742), .A2(new_n374), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1065), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n726), .B1(new_n1072), .B2(new_n728), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1055), .B(new_n1073), .C1(new_n352), .C2(new_n816), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1054), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1044), .A2(new_n1052), .A3(new_n1047), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1052), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT118), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT118), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1051), .A2(new_n1079), .A3(new_n1053), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT116), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1049), .A2(new_n865), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1038), .B1(new_n1082), .B2(new_n1050), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1049), .A2(new_n865), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1052), .A2(new_n1046), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n870), .A2(new_n635), .A3(new_n885), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1081), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g0889(.A(KEYINPUT116), .B(new_n1087), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1078), .A2(new_n1080), .A3(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT119), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1051), .B(new_n1053), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT117), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n688), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1094), .B2(new_n688), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1075), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(KEYINPUT121), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n884), .A2(new_n867), .A3(new_n868), .A4(new_n861), .ZN(new_n1102));
  INV_X1    g0902(.A(G330), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n877), .B2(new_n879), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n869), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n437), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n634), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n414), .A2(new_n844), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT55), .Z(new_n1109));
  XNOR2_X1  g0909(.A(new_n1107), .B(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1102), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1101), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1112), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1104), .A2(new_n869), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1104), .A2(new_n869), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1102), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(KEYINPUT121), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n1088), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT122), .B1(new_n1094), .B2(new_n1088), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n689), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(KEYINPUT57), .B1(new_n1113), .B2(new_n1114), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n947), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1112), .A2(new_n788), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n963), .B1(new_n355), .B2(new_n768), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n996), .C1(new_n889), .C2(new_n752), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n957), .A2(G58), .ZN(new_n1134));
  AOI21_X1  g0934(.A(G41), .B1(new_n764), .B2(G107), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n754), .C2(new_n374), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n735), .A2(new_n778), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n1133), .A2(new_n283), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT58), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n260), .B1(new_n276), .B2(new_n278), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n223), .B1(new_n1140), .B2(G41), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n757), .A2(G150), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n802), .A2(new_n1059), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n768), .A2(G137), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n753), .A2(G132), .B1(G128), .B2(new_n764), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G125), .B2(new_n751), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT59), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G33), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G41), .B1(new_n810), .B2(G124), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n736), .C2(new_n760), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n728), .B1(new_n1139), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n815), .A2(new_n201), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1131), .A2(new_n725), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1130), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1129), .A2(new_n1158), .ZN(G375));
  AOI211_X1 g0959(.A(new_n964), .B(new_n992), .C1(new_n461), .C2(new_n753), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n802), .A2(G97), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n810), .A2(G303), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n264), .B1(new_n741), .B2(new_n778), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n751), .B2(G294), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n742), .A2(new_n364), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n752), .A2(new_n804), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1134), .B1(new_n409), .B2(new_n742), .C1(new_n754), .C2(new_n1060), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G50), .B2(new_n757), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n810), .A2(G128), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n802), .A2(G159), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n280), .B1(G137), .B2(new_n764), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1165), .A2(new_n1166), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n726), .B1(new_n1174), .B2(new_n728), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(G68), .B2(new_n816), .C1(new_n1039), .C2(new_n789), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1086), .B2(new_n947), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1083), .A2(new_n1087), .A3(new_n1085), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1091), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n927), .B(KEYINPUT123), .Z(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(G381));
  AOI21_X1  g0982(.A(new_n1157), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1099), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1186));
  OR2_X1    g0986(.A1(G393), .A2(G396), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(G407));
  NOR2_X1   g0989(.A1(new_n662), .A2(G343), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(KEYINPUT124), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT124), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1184), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(G407), .A2(new_n1191), .A3(G213), .A4(new_n1194), .ZN(G409));
  AOI21_X1  g0995(.A(new_n1033), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1094), .A2(new_n1088), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n1088), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1199), .A2(new_n1200), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1181), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1196), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1099), .A3(new_n1156), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1193), .C1(new_n1183), .C2(new_n1099), .ZN(new_n1205));
  XOR2_X1   g1005(.A(G384), .B(KEYINPUT125), .Z(new_n1206));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1179), .A2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n689), .B(new_n1208), .C1(new_n1180), .C2(KEYINPUT60), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1178), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1206), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1180), .B2(KEYINPUT60), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n688), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1178), .A3(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1190), .A2(G2897), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1211), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1205), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT63), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1190), .B1(G375), .B2(G378), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1204), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G390), .A2(new_n948), .A3(new_n977), .ZN(new_n1227));
  INV_X1    g1027(.A(G396), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(G393), .B(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(G387), .A2(new_n1035), .A3(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G387), .A2(new_n1035), .B1(new_n1229), .B2(KEYINPUT126), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(KEYINPUT126), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1222), .A2(KEYINPUT63), .A3(new_n1204), .A4(new_n1223), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1225), .A2(new_n1226), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1222), .A2(new_n1238), .A3(new_n1204), .A4(new_n1223), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1223), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT62), .B1(new_n1205), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT127), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT127), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1244), .B(KEYINPUT61), .C1(new_n1205), .C2(new_n1219), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1237), .B1(new_n1246), .B2(new_n1235), .ZN(G405));
  NAND2_X1  g1047(.A1(G375), .A2(G378), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1235), .A2(new_n1184), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1184), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(new_n1240), .ZN(G402));
endmodule


