//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT24), .A3(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n205), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n208), .A2(new_n216), .A3(KEYINPUT25), .A4(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(new_n217), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n224), .B2(new_n215), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n205), .B(KEYINPUT65), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n218), .B(new_n227), .C1(new_n228), .C2(KEYINPUT26), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT27), .B(G183gat), .Z(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n233));
  AOI21_X1  g032(.A(G190gat), .B1(new_n233), .B2(KEYINPUT66), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT28), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n230), .A2(new_n236), .A3(G190gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n229), .B(new_n212), .C1(new_n235), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(KEYINPUT67), .B2(KEYINPUT1), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n241), .B(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n238), .B2(new_n226), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT34), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n249), .B2(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n245), .A2(new_n249), .A3(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT32), .ZN(new_n255));
  INV_X1    g054(.A(new_n252), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n249), .B(new_n256), .C1(new_n245), .C2(new_n247), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n248), .B2(new_n249), .ZN(new_n259));
  INV_X1    g058(.A(new_n257), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT32), .B(new_n254), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n258), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(new_n258), .B2(new_n261), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n203), .B(new_n204), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n258), .A2(new_n261), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n267), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n261), .A3(new_n268), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(KEYINPUT69), .A3(new_n202), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT80), .B(G50gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G155gat), .B(G162gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n283), .A2(KEYINPUT73), .B1(KEYINPUT2), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G141gat), .B(G148gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n287), .C1(KEYINPUT73), .C2(new_n283), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  INV_X1    g090(.A(new_n283), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n286), .B2(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n289), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT81), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n302), .A2(new_n304), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n291), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n315), .A3(new_n307), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G228gat), .ZN(new_n318));
  INV_X1    g117(.A(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n291), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n310), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n297), .A2(new_n307), .B1(new_n323), .B2(new_n310), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT82), .A3(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n322), .A2(new_n330), .A3(G22gat), .ZN(new_n331));
  INV_X1    g130(.A(G22gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n325), .A2(new_n326), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT82), .B1(new_n328), .B2(new_n320), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n321), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n282), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(G22gat), .B1(new_n322), .B2(new_n330), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n332), .A3(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .A4(new_n281), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(KEYINPUT83), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n310), .A2(new_n246), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n290), .A2(new_n244), .A3(new_n293), .A4(new_n294), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n350), .B(KEYINPUT75), .Z(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(KEYINPUT76), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n246), .A3(new_n295), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n355), .A2(new_n356), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n358), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n363), .A2(KEYINPUT5), .A3(new_n351), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365));
  INV_X1    g164(.A(new_n354), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n359), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n354), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n352), .A2(new_n362), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G85gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  AOI21_X1  g173(.A(new_n345), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n364), .A2(new_n369), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n358), .A3(new_n356), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n366), .A2(new_n359), .A3(new_n360), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n352), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n376), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI211_X1 g182(.A(KEYINPUT84), .B(new_n374), .C1(new_n377), .C2(new_n380), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n375), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n345), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  INV_X1    g186(.A(G64gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G92gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT72), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n239), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n307), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n226), .B2(new_n238), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT37), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(KEYINPUT37), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT38), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n404), .A2(new_n405), .B1(new_n392), .B2(new_n401), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n385), .A2(new_n386), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT39), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n351), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n347), .A2(new_n356), .A3(new_n348), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT39), .B(new_n413), .C1(new_n409), .C2(new_n356), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n415), .A2(KEYINPUT40), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n412), .A2(new_n414), .A3(new_n374), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT84), .B1(new_n370), .B2(new_n374), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n381), .A2(new_n376), .A3(new_n382), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n409), .A2(new_n356), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n382), .B1(new_n423), .B2(new_n411), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n424), .A2(new_n415), .A3(KEYINPUT40), .A4(new_n414), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT30), .B1(new_n401), .B2(new_n392), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n392), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n419), .A2(new_n422), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n276), .B(new_n344), .C1(new_n408), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n375), .B1(new_n374), .B2(new_n370), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n386), .ZN(new_n432));
  INV_X1    g231(.A(new_n428), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n344), .A2(new_n275), .A3(new_n271), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n339), .A2(new_n340), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(new_n282), .B1(KEYINPUT83), .B2(new_n331), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n269), .A2(new_n270), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(KEYINPUT35), .A3(new_n342), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n438), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n344), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n428), .B1(new_n385), .B2(new_n386), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT35), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n430), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(KEYINPUT86), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(KEYINPUT86), .ZN(new_n449));
  NOR3_X1   g248(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G29gat), .ZN(new_n452));
  INV_X1    g251(.A(G36gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT15), .B(new_n446), .C1(new_n451), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n446), .A2(new_n459), .A3(KEYINPUT15), .ZN(new_n460));
  OR3_X1    g259(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n454), .B1(new_n461), .B2(new_n447), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n457), .A2(new_n458), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT17), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT88), .B(new_n467), .C1(new_n455), .C2(new_n463), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(G1gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT90), .ZN(new_n473));
  INV_X1    g272(.A(G8gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n475), .A3(new_n471), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n469), .A2(G1gat), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(KEYINPUT89), .B2(G8gat), .ZN(new_n479));
  AND4_X1   g278(.A1(KEYINPUT89), .A2(new_n478), .A3(G8gat), .A4(new_n472), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n466), .A2(new_n468), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT18), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n482), .B(new_n464), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n484), .B(KEYINPUT13), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n481), .A2(KEYINPUT18), .A3(new_n483), .A4(new_n484), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT11), .B(G169gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G197gat), .ZN(new_n495));
  XOR2_X1   g294(.A(G113gat), .B(G141gat), .Z(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT12), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n487), .A2(new_n498), .A3(new_n491), .A4(new_n492), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT91), .B1(new_n445), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n435), .A2(new_n439), .ZN(new_n505));
  INV_X1    g304(.A(new_n434), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n442), .A2(new_n443), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n408), .A2(new_n429), .ZN(new_n511));
  INV_X1    g310(.A(new_n344), .ZN(new_n512));
  INV_X1    g311(.A(new_n276), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n507), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n502), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n504), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT95), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(G85gat), .A3(G92gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  INV_X1    g323(.A(G85gat), .ZN(new_n525));
  AOI22_X1  g324(.A1(KEYINPUT8), .A2(new_n524), .B1(new_n525), .B2(new_n390), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(KEYINPUT95), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n524), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n523), .A2(new_n532), .A3(new_n526), .A4(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n466), .B2(new_n468), .ZN(new_n535));
  XOR2_X1   g334(.A(G190gat), .B(G218gat), .Z(new_n536));
  INV_X1    g335(.A(new_n534), .ZN(new_n537));
  AND2_X1   g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n464), .A2(new_n537), .B1(KEYINPUT41), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n536), .B1(new_n535), .B2(new_n539), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI211_X1 g345(.A(KEYINPUT97), .B(new_n536), .C1(new_n535), .C2(new_n539), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n542), .A2(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n538), .A2(KEYINPUT41), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI221_X1 g352(.A(new_n551), .B1(new_n546), .B2(new_n547), .C1(new_n542), .C2(new_n543), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n556));
  INV_X1    g355(.A(G57gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(G64gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n388), .A2(G57gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n388), .A2(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n561), .A2(new_n562), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n565), .A2(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT21), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(G183gat), .B1(new_n482), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT19), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n209), .B(new_n574), .C1(new_n479), .C2(new_n480), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n556), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n573), .A2(KEYINPUT21), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n582), .B2(new_n584), .ZN(new_n588));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT94), .B(G211gat), .Z(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n590), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n587), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT20), .B1(new_n583), .B2(new_n579), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n580), .A2(new_n581), .A3(new_n556), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n585), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n555), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n595), .B1(new_n587), .B2(new_n588), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n600), .A3(new_n594), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n555), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n537), .A2(KEYINPUT10), .A3(new_n573), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n565), .A2(new_n569), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n533), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n571), .A2(new_n572), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n534), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n573), .A2(KEYINPUT99), .A3(new_n533), .A4(new_n531), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n617), .A2(new_n619), .A3(new_n622), .A4(new_n618), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n611), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n617), .A2(new_n619), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT101), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G120gat), .ZN(new_n634));
  INV_X1    g433(.A(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n628), .A2(new_n630), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n609), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n518), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n432), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n433), .ZN(new_n647));
  NAND2_X1  g446(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n470), .A2(new_n474), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n647), .A2(KEYINPUT42), .A3(new_n648), .A4(new_n649), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n652), .B(new_n653), .C1(new_n474), .C2(new_n647), .ZN(G1325gat));
  AOI21_X1  g453(.A(G15gat), .B1(new_n643), .B2(new_n438), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n642), .A2(new_n513), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(G15gat), .B2(new_n656), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n512), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n607), .A2(new_n640), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n504), .B2(new_n517), .ZN(new_n664));
  INV_X1    g463(.A(new_n555), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n452), .A3(new_n644), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n661), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n667), .A3(KEYINPUT45), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n445), .B2(new_n555), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n515), .A2(KEYINPUT44), .A3(new_n665), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n662), .A2(new_n502), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679), .B2(new_n432), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n670), .A2(new_n672), .A3(new_n680), .ZN(G1328gat));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n665), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(G36gat), .A3(new_n433), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n679), .B2(new_n433), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(G1329gat));
  OR3_X1    g487(.A1(new_n682), .A2(G43gat), .A3(new_n441), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690));
  OAI21_X1  g489(.A(G43gat), .B1(new_n679), .B2(new_n513), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(G1330gat));
  NAND4_X1  g493(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n344), .A4(new_n678), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n674), .A2(new_n344), .A3(new_n675), .A4(new_n678), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(G50gat), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n512), .A2(G50gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n664), .A2(new_n665), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(KEYINPUT48), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n696), .A2(G50gat), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT48), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n701), .A4(KEYINPUT48), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n609), .A2(new_n502), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n515), .A2(new_n640), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n432), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n557), .ZN(G1332gat));
  AOI211_X1 g512(.A(new_n433), .B(new_n711), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n711), .B2(new_n513), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n711), .A2(G71gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n441), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g519(.A1(new_n711), .A2(new_n512), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(G78gat), .Z(G1335gat));
  AND3_X1   g521(.A1(new_n674), .A2(new_n640), .A3(new_n675), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n607), .A2(new_n502), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n644), .A4(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n674), .A2(new_n640), .A3(new_n675), .A4(new_n724), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n432), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(G85gat), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n515), .A2(new_n665), .A3(new_n724), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT51), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n515), .A2(new_n732), .A3(new_n665), .A4(new_n724), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n640), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n525), .A3(new_n644), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n735), .ZN(G1336gat));
  NOR2_X1   g535(.A1(new_n433), .A2(G92gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n731), .A2(new_n640), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n740));
  OAI21_X1  g539(.A(G92gat), .B1(new_n727), .B2(new_n433), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n741), .A2(new_n742), .A3(new_n738), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n738), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n738), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n747));
  INV_X1    g546(.A(new_n740), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n741), .A2(new_n742), .A3(new_n738), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n745), .A2(new_n750), .ZN(G1337gat));
  INV_X1    g550(.A(G99gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n752), .A3(new_n438), .ZN(new_n753));
  OAI21_X1  g552(.A(G99gat), .B1(new_n727), .B2(new_n513), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1338gat));
  NOR2_X1   g554(.A1(new_n512), .A2(G106gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G106gat), .B1(new_n727), .B2(new_n512), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT53), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n723), .A2(KEYINPUT109), .A3(new_n344), .A4(new_n724), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n727), .B2(new_n512), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(G106gat), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT53), .B1(new_n734), .B2(new_n756), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n767), .B2(new_n768), .ZN(G1339gat));
  INV_X1    g568(.A(new_n639), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n625), .B(new_n611), .C1(new_n621), .C2(new_n623), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n627), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n624), .A2(KEYINPUT54), .A3(new_n626), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT111), .B1(new_n774), .B2(new_n636), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n621), .A2(new_n623), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n610), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n772), .A3(new_n625), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n637), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n773), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n770), .B1(new_n781), .B2(KEYINPUT55), .ZN(new_n782));
  INV_X1    g581(.A(new_n773), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n636), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n778), .B2(new_n637), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(new_n788), .A3(new_n502), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n488), .A2(new_n490), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n484), .B1(new_n481), .B2(new_n483), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n497), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n501), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n640), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n665), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n665), .A2(new_n782), .A3(new_n788), .A4(new_n793), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n607), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n640), .A2(new_n793), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n502), .B1(new_n781), .B2(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n801), .B1(new_n803), .B2(new_n782), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n800), .B(new_n796), .C1(new_n804), .C2(new_n665), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n798), .A2(new_n799), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n640), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n604), .A2(new_n503), .A3(new_n608), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n442), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n644), .A2(new_n433), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n502), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n640), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n607), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT113), .A2(G127gat), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n818), .B(new_n819), .Z(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n810), .A2(new_n821), .A3(new_n665), .A4(new_n812), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n810), .A2(new_n665), .A3(new_n812), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT114), .B1(new_n825), .B2(G134gat), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n825), .A2(KEYINPUT114), .A3(G134gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n824), .B(KEYINPUT115), .C1(new_n826), .C2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1343gat));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n835), .A3(new_n344), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n811), .A2(new_n276), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n639), .B1(new_n786), .B2(new_n787), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n794), .B1(new_n839), .B2(new_n802), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n555), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n607), .B1(new_n841), .B2(new_n796), .ZN(new_n842));
  INV_X1    g641(.A(new_n808), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n344), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n838), .B1(new_n844), .B2(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n502), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G141gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n834), .A2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n512), .B1(new_n806), .B2(new_n808), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n503), .A2(G141gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n837), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n809), .A2(new_n344), .A3(new_n837), .A4(new_n852), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n847), .A2(new_n849), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n846), .A2(new_n857), .A3(G141gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n834), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n848), .B1(new_n846), .B2(G141gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n833), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n858), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n855), .A2(new_n853), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n861), .C1(new_n866), .C2(new_n834), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n809), .A2(new_n344), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n838), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n635), .A3(new_n640), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n842), .B2(new_n843), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n799), .B1(new_n795), .B2(new_n797), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT119), .A3(new_n808), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(KEYINPUT57), .A2(new_n869), .B1(new_n877), .B2(new_n344), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n640), .A3(new_n837), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n836), .A2(new_n845), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n635), .C1(new_n881), .C2(new_n640), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n880), .B2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(G155gat), .B1(new_n870), .B2(new_n607), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n607), .A2(G155gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n870), .B2(new_n665), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n665), .A2(G162gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n881), .B2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n644), .A2(new_n433), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n810), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G169gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n502), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n890), .B(KEYINPUT120), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n810), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n503), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n891), .B2(new_n640), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n807), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(G176gat), .B2(new_n899), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n799), .A2(new_n230), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G183gat), .B1(new_n895), .B2(new_n799), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n906));
  NAND2_X1  g705(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n907), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n903), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n908), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n210), .A3(new_n665), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT123), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n917));
  OAI211_X1 g716(.A(G190gat), .B(new_n917), .C1(new_n895), .C2(new_n555), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n877), .A2(new_n344), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n894), .A2(new_n513), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n503), .ZN(new_n927));
  AND4_X1   g726(.A1(new_n344), .A2(new_n809), .A3(new_n513), .A4(new_n890), .ZN(new_n928));
  INV_X1    g727(.A(G197gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n502), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(new_n640), .ZN(new_n933));
  AND2_X1   g732(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n934));
  NOR2_X1   g733(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n878), .A2(new_n640), .A3(new_n925), .ZN(new_n937));
  OAI221_X1 g736(.A(new_n936), .B1(new_n934), .B2(new_n933), .C1(new_n937), .C2(new_n932), .ZN(G1353gat));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n939), .A3(new_n607), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n926), .B2(new_n799), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n878), .A2(KEYINPUT126), .A3(new_n607), .A4(new_n925), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(G211gat), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n928), .B2(new_n665), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT127), .Z(new_n950));
  INV_X1    g749(.A(new_n926), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n665), .A2(G218gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1355gat));
endmodule


