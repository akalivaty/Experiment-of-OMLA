//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT73), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G237), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT73), .ZN(new_n193));
  OAI211_X1 g007(.A(G214), .B(new_n189), .C1(new_n191), .C2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(KEYINPUT73), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G237), .ZN(new_n198));
  AOI21_X1  g012(.A(G953), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(G143), .B1(new_n199), .B2(G214), .ZN(new_n200));
  OAI21_X1  g014(.A(G131), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(G143), .A3(G214), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(KEYINPUT77), .A3(G125), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT16), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n207), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT19), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(KEYINPUT92), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n213), .A2(new_n214), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n207), .B(new_n222), .C1(new_n224), .C2(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n206), .A2(new_n219), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n202), .A2(new_n204), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT18), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AOI211_X1 g045(.A(KEYINPUT88), .B(new_n229), .C1(new_n202), .C2(new_n204), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n213), .A2(G146), .A3(new_n214), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n220), .B2(new_n207), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n213), .A2(new_n234), .A3(G146), .A4(new_n214), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n236), .A2(KEYINPUT90), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT90), .B1(new_n236), .B2(new_n237), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n231), .A2(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n202), .A2(new_n204), .A3(new_n229), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT91), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT91), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n202), .A2(new_n243), .A3(new_n204), .A4(new_n229), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n226), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G113), .B(G122), .ZN(new_n247));
  INV_X1    g061(.A(G104), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n201), .A2(new_n252), .A3(new_n205), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n215), .A2(new_n207), .A3(new_n217), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n218), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n228), .A2(KEYINPUT17), .A3(G131), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(new_n249), .C1(new_n240), .C2(new_n245), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n188), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT93), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n230), .B1(new_n196), .B2(new_n200), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT88), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n228), .A2(new_n227), .A3(new_n230), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n242), .A2(new_n244), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n236), .A2(new_n237), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n236), .A2(KEYINPUT90), .A3(new_n237), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n249), .B1(new_n274), .B2(new_n226), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n187), .B1(new_n263), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT20), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n261), .B(new_n187), .C1(new_n263), .C2(new_n275), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n262), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n249), .B1(new_n274), .B2(new_n258), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n263), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G475), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G116), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n287), .B2(G116), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT96), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G122), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT96), .B1(new_n293), .B2(KEYINPUT14), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT97), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n290), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(KEYINPUT96), .A3(KEYINPUT14), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n288), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n293), .A2(KEYINPUT14), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G107), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n195), .A2(G128), .ZN(new_n303));
  INV_X1    g117(.A(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G134), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G107), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n288), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT13), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n303), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n195), .A2(KEYINPUT13), .A3(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n305), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT94), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n322), .A3(G134), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n303), .A2(new_n305), .A3(new_n325), .A4(new_n308), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n293), .A2(new_n288), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n312), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n309), .A2(KEYINPUT95), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n326), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT9), .B(G234), .ZN(new_n332));
  INV_X1    g146(.A(G217), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n332), .A2(new_n333), .A3(G953), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n313), .B1(new_n301), .B2(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n326), .A3(new_n330), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n321), .B2(new_n323), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n281), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n343), .A2(KEYINPUT15), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  AND2_X1   g159(.A1(new_n189), .A2(G952), .ZN(new_n346));
  NAND2_X1  g160(.A1(G234), .A2(G237), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(G902), .A3(G953), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT21), .B(G898), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n286), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G221), .ZN(new_n356));
  INV_X1    g170(.A(new_n332), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n281), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n281), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G140), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n189), .A2(G227), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT12), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n207), .A2(G143), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT69), .B1(new_n367), .B2(KEYINPUT1), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT69), .B(KEYINPUT1), .C1(new_n195), .C2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G128), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n207), .B2(G143), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n195), .A2(KEYINPUT66), .A3(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT65), .B1(new_n195), .B2(G146), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT65), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n207), .A3(G143), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n304), .A2(KEYINPUT1), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n379), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(new_n248), .B2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n311), .A3(G104), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n248), .A2(G107), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n248), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n311), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n374), .A2(new_n383), .A3(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n195), .A2(KEYINPUT66), .A3(G146), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT66), .B1(new_n195), .B2(G146), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n379), .B(new_n381), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n367), .A2(KEYINPUT1), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(KEYINPUT84), .A3(new_n399), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n383), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n393), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n394), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT11), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n308), .B2(G137), .ZN(new_n408));
  AOI21_X1  g222(.A(G131), .B1(new_n308), .B2(G137), .ZN(new_n409));
  INV_X1    g223(.A(G137), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT11), .A3(G134), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT68), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n308), .A2(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G131), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n366), .B1(new_n406), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n397), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n400), .A2(new_n401), .B1(new_n423), .B2(new_n382), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n393), .B1(new_n424), .B2(new_n403), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT12), .B(new_n420), .C1(new_n425), .C2(new_n394), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n379), .A2(new_n381), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n428), .A2(new_n378), .B1(G128), .B2(new_n398), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n383), .B1(new_n429), .B2(KEYINPUT84), .ZN(new_n430));
  INV_X1    g244(.A(new_n403), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n405), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G101), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(new_n439), .A3(new_n436), .A4(G101), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n435), .B2(G101), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n438), .A2(new_n440), .B1(new_n389), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n195), .A2(G146), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n207), .B2(G143), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(KEYINPUT0), .A2(G128), .ZN(new_n448));
  NOR2_X1   g262(.A1(KEYINPUT0), .A2(G128), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n378), .A2(new_n448), .A3(new_n379), .A4(new_n381), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT67), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n428), .A2(new_n453), .A3(new_n448), .A4(new_n378), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n373), .A2(new_n371), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n383), .B1(new_n456), .B2(new_n447), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n393), .A2(new_n433), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n442), .A2(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n434), .A2(new_n421), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n365), .B1(new_n427), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT82), .B1(new_n427), .B2(new_n460), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n455), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT10), .B1(new_n404), .B2(new_n405), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n465), .A2(new_n466), .A3(new_n420), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n421), .B1(new_n434), .B2(new_n459), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n364), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n364), .A2(new_n461), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n360), .B1(new_n470), .B2(G469), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n427), .A2(KEYINPUT85), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT85), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n422), .A2(new_n426), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n460), .A2(new_n364), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n420), .B1(new_n465), .B2(new_n466), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n364), .B1(new_n477), .B2(new_n460), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n359), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n358), .B1(new_n471), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n438), .A2(new_n440), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT2), .B(G113), .Z(new_n486));
  XNOR2_X1  g300(.A(G116), .B(G119), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n441), .A2(new_n389), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g305(.A(G119), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G116), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n491), .B(G113), .C1(KEYINPUT5), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n486), .A2(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n405), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G122), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n405), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n494), .B(new_n495), .C1(KEYINPUT86), .C2(new_n393), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n497), .B(KEYINPUT8), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n374), .A2(new_n210), .A3(new_n383), .ZN(new_n505));
  INV_X1    g319(.A(G224), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(G953), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n505), .B(new_n509), .C1(new_n455), .C2(new_n210), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n498), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n505), .A2(KEYINPUT87), .B1(new_n508), .B2(new_n507), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n455), .B2(new_n210), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n490), .A2(new_n496), .ZN(new_n518));
  INV_X1    g332(.A(new_n497), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n514), .A2(new_n507), .ZN(new_n524));
  OAI221_X1 g338(.A(new_n505), .B1(new_n506), .B2(G953), .C1(new_n455), .C2(new_n210), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G210), .B1(G237), .B2(G902), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n517), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n517), .B2(new_n527), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n484), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n355), .A2(new_n483), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n452), .A2(new_n454), .ZN(new_n534));
  INV_X1    g348(.A(new_n450), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n420), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n488), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n410), .A2(G134), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n203), .B1(new_n539), .B2(new_n417), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n414), .B2(new_n415), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n457), .B1(new_n541), .B2(KEYINPUT70), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n543), .B(new_n540), .C1(new_n414), .C2(new_n415), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT72), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n540), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n416), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n543), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(KEYINPUT70), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n457), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n488), .B1(new_n455), .B2(new_n420), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n199), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT27), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT26), .B(G101), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n546), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n457), .A2(new_n541), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n536), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n537), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n455), .B2(new_n420), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n551), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n551), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT31), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n455), .A2(new_n420), .B1(new_n457), .B2(new_n541), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n488), .B1(new_n571), .B2(KEYINPUT30), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT71), .B1(new_n573), .B2(new_n545), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n551), .A2(new_n565), .A3(new_n564), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n546), .A2(new_n554), .A3(new_n558), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT31), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT28), .B1(new_n551), .B2(new_n552), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n488), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n546), .A2(new_n580), .A3(new_n554), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n581), .B2(KEYINPUT28), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n570), .B(new_n578), .C1(new_n582), .C2(new_n558), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n534), .A2(new_n420), .A3(new_n535), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n488), .B1(new_n545), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n546), .A2(new_n554), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n579), .B1(new_n591), .B2(KEYINPUT28), .ZN(new_n592));
  INV_X1    g406(.A(new_n558), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n546), .A2(new_n554), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n593), .B1(new_n576), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n594), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n579), .B(new_n593), .C1(new_n581), .C2(KEYINPUT28), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n583), .A2(KEYINPUT32), .A3(new_n584), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n588), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT22), .B(G137), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n220), .A2(new_n207), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n304), .A2(G119), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n492), .A2(G128), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G110), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT24), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G110), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT75), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT75), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n616), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n614), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT23), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n492), .B2(G128), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n304), .A2(KEYINPUT23), .A3(G119), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n612), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(G110), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n610), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT78), .B1(new_n629), .B2(new_n218), .ZN(new_n630));
  INV_X1    g444(.A(new_n610), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n627), .A2(G110), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n616), .A2(new_n618), .A3(new_n621), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n621), .B1(new_n616), .B2(new_n618), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n613), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT78), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n219), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(G110), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT76), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n633), .A2(new_n634), .A3(new_n613), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT76), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n627), .B2(G110), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n218), .B2(new_n255), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n609), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n629), .A2(KEYINPUT78), .A3(new_n218), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n637), .B1(new_n636), .B2(new_n219), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT79), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT79), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n639), .A2(new_n652), .A3(new_n646), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n647), .B1(new_n654), .B2(new_n609), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n333), .B1(G234), .B2(new_n281), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(G902), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n605), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n608), .B1(new_n651), .B2(new_n653), .ZN(new_n660));
  OAI211_X1 g474(.A(KEYINPUT80), .B(new_n657), .C1(new_n660), .C2(new_n647), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n650), .A2(KEYINPUT79), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n652), .B1(new_n639), .B2(new_n646), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n609), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n647), .ZN(new_n666));
  AOI21_X1  g480(.A(G902), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT25), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n656), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n281), .B1(new_n660), .B2(new_n647), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(KEYINPUT25), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n662), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n604), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(KEYINPUT81), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT81), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n604), .B2(new_n673), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n533), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT98), .B(G101), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G3));
  NAND2_X1  g494(.A1(new_n570), .A2(new_n578), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n581), .A2(KEYINPUT28), .ZN(new_n682));
  INV_X1    g496(.A(new_n579), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n558), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n281), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n685), .A2(G472), .B1(new_n584), .B2(new_n583), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n482), .A2(new_n673), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n484), .ZN(new_n688));
  INV_X1    g502(.A(new_n528), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n690));
  INV_X1    g504(.A(new_n516), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n498), .A2(new_n504), .A3(new_n510), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n281), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n688), .B1(new_n694), .B2(new_n529), .ZN(new_n695));
  INV_X1    g509(.A(new_n353), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n700));
  AOI21_X1  g514(.A(new_n334), .B1(new_n315), .B2(new_n331), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n337), .A2(new_n339), .A3(new_n336), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n335), .A2(new_n340), .A3(KEYINPUT33), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n699), .B1(new_n341), .B2(new_n700), .ZN(new_n706));
  OAI21_X1  g520(.A(G478), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n342), .A2(G478), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n343), .A2(new_n281), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n285), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n687), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT34), .B(G104), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G6));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n279), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n260), .A2(KEYINPUT101), .A3(new_n261), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n262), .A2(new_n718), .A3(new_n278), .A4(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n284), .A3(new_n345), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n687), .A2(new_n697), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT35), .B(G107), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G9));
  NAND3_X1  g538(.A1(new_n482), .A2(new_n686), .A3(new_n695), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n654), .A2(KEYINPUT36), .A3(new_n609), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n609), .A2(KEYINPUT36), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n651), .B2(new_n653), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n657), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n656), .B1(new_n667), .B2(new_n668), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n671), .A2(KEYINPUT25), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n286), .A2(new_n354), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n725), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT37), .B(G110), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G12));
  XOR2_X1   g550(.A(KEYINPUT102), .B(G900), .Z(new_n737));
  AOI21_X1  g551(.A(new_n349), .B1(new_n351), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n284), .A2(new_n720), .A3(new_n345), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n672), .A2(new_n669), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n532), .B1(new_n741), .B2(new_n729), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n604), .A2(new_n740), .A3(new_n482), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G128), .ZN(G30));
  XOR2_X1   g558(.A(new_n738), .B(KEYINPUT39), .Z(new_n745));
  NAND2_X1  g559(.A1(new_n482), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT40), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n746), .B(KEYINPUT104), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT40), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n576), .A2(new_n597), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n593), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n281), .B1(new_n591), .B2(new_n558), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n588), .A2(new_n603), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT103), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n530), .A2(new_n531), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT38), .Z(new_n761));
  INV_X1    g575(.A(new_n345), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n286), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n732), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n763), .A3(new_n484), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n750), .A2(new_n752), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G143), .ZN(G45));
  AOI211_X1 g582(.A(new_n738), .B(new_n711), .C1(new_n280), .C2(new_n284), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n604), .A2(new_n769), .A3(new_n482), .A4(new_n742), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G146), .ZN(G48));
  AOI21_X1  g585(.A(new_n358), .B1(new_n480), .B2(new_n359), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n480), .B2(KEYINPUT105), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n473), .B1(new_n422), .B2(new_n426), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n460), .A2(new_n364), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n478), .B1(new_n776), .B2(new_n474), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT105), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(G902), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT106), .B(new_n772), .C1(new_n773), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n480), .A2(KEYINPUT105), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n778), .B1(new_n777), .B2(G902), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(G469), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT106), .B1(new_n784), .B2(new_n772), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT107), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n674), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n772), .B1(new_n773), .B2(new_n779), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n780), .ZN(new_n792));
  INV_X1    g606(.A(new_n713), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n786), .A2(new_n787), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT41), .B(G113), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G15));
  NAND2_X1  g610(.A1(new_n786), .A2(new_n792), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n721), .A2(new_n697), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n604), .A3(new_n673), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G116), .ZN(G18));
  NOR3_X1   g616(.A1(new_n781), .A2(new_n785), .A3(new_n532), .ZN(new_n803));
  INV_X1    g617(.A(new_n733), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n604), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G119), .ZN(G21));
  NOR2_X1   g620(.A1(new_n592), .A2(new_n558), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n584), .B1(new_n681), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT108), .B1(new_n685), .B2(G472), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(G472), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n810), .B(new_n811), .C1(new_n583), .C2(new_n281), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n673), .B(new_n808), .C1(new_n809), .C2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n285), .A2(new_n695), .A3(new_n696), .A4(new_n345), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n798), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G122), .ZN(G24));
  NAND2_X1  g631(.A1(new_n685), .A2(G472), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n810), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n685), .A2(KEYINPUT108), .A3(G472), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n732), .A3(new_n769), .A4(new_n808), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n790), .A2(new_n695), .A3(new_n780), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n210), .ZN(G27));
  INV_X1    g639(.A(KEYINPUT42), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n694), .A2(new_n484), .A3(new_n529), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n694), .A2(new_n829), .A3(new_n529), .A4(new_n484), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n604), .A2(new_n831), .A3(new_n673), .A4(new_n482), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n285), .A2(new_n712), .A3(new_n739), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT32), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n585), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n602), .A3(new_n603), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n673), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n828), .A2(new_n830), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n483), .A2(new_n826), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G131), .ZN(G33));
  AND4_X1   g658(.A1(new_n604), .A2(new_n831), .A3(new_n673), .A4(new_n482), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n740), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G134), .ZN(G36));
  OR2_X1    g661(.A1(new_n285), .A2(KEYINPUT111), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT43), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n286), .A2(new_n712), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n764), .A2(new_n686), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT44), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n839), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n470), .A2(KEYINPUT45), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n359), .B1(new_n470), .B2(KEYINPUT45), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n360), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n481), .B1(new_n858), .B2(KEYINPUT46), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(KEYINPUT46), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT110), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT110), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n358), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n745), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n850), .A2(new_n851), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n848), .A2(new_n849), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n286), .B2(new_n712), .ZN(new_n869));
  OAI211_X1 g683(.A(KEYINPUT44), .B(new_n853), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n855), .B(new_n866), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(G137), .ZN(G39));
  NAND3_X1  g689(.A1(new_n864), .A2(KEYINPUT47), .A3(new_n865), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT47), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n863), .B2(new_n358), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n588), .A2(new_n602), .A3(new_n603), .ZN(new_n880));
  INV_X1    g694(.A(new_n673), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n840), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(G140), .ZN(G42));
  NOR2_X1   g697(.A1(new_n781), .A2(new_n785), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n831), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT118), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n348), .B1(new_n885), .B2(KEYINPUT118), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n852), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n732), .B(new_n808), .C1(new_n809), .C2(new_n812), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n850), .A2(new_n851), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n868), .A2(new_n286), .A3(new_n712), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n348), .B(new_n813), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n761), .A2(new_n484), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n884), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT50), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n673), .A2(new_n886), .A3(new_n759), .A4(new_n887), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n285), .A2(new_n712), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n784), .A2(new_n481), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n876), .B(new_n878), .C1(new_n865), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n831), .A3(new_n898), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n895), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n895), .A2(new_n906), .A3(KEYINPUT51), .A4(new_n909), .ZN(new_n913));
  INV_X1    g727(.A(new_n838), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n890), .B2(new_n891), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT48), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n904), .A2(new_n285), .A3(new_n712), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n898), .A2(new_n803), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n346), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n915), .B2(KEYINPUT48), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n912), .A2(new_n913), .A3(new_n916), .A4(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n786), .B(new_n792), .C1(new_n815), .C2(new_n800), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n843), .A3(new_n794), .A4(new_n805), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n280), .A2(new_n284), .A3(new_n345), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n926), .B2(new_n698), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n697), .A3(KEYINPUT115), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n687), .A3(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n713), .A2(new_n687), .B1(new_n725), .B2(new_n733), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n345), .A2(new_n738), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n732), .A2(new_n284), .A3(new_n720), .A4(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n880), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n483), .A2(new_n839), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n845), .A2(new_n740), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n893), .A2(new_n833), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n935), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n931), .A2(new_n936), .A3(new_n678), .A4(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n923), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT52), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n803), .A2(new_n937), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n285), .A2(new_n695), .A3(new_n345), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n732), .A2(new_n738), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n757), .A3(new_n944), .A4(new_n482), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n945), .A2(new_n743), .A3(new_n770), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n743), .A3(new_n770), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n824), .A2(new_n948), .A3(KEYINPUT52), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT116), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n942), .A2(new_n946), .A3(new_n941), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT52), .B1(new_n824), .B2(new_n948), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT116), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n940), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT53), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT53), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n947), .A2(new_n949), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n940), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(KEYINPUT54), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n955), .A2(new_n957), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n923), .A2(KEYINPUT117), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n939), .A2(new_n957), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n923), .A2(KEYINPUT117), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n958), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  OAI22_X1  g782(.A1(new_n921), .A2(new_n968), .B1(G952), .B2(G953), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n673), .A2(new_n865), .A3(new_n484), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT113), .Z(new_n971));
  AOI21_X1  g785(.A(new_n851), .B1(new_n907), .B2(KEYINPUT49), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT114), .Z(new_n974));
  INV_X1    g788(.A(new_n761), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n907), .A2(KEYINPUT49), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n974), .A2(new_n759), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n969), .A2(new_n977), .ZN(G75));
  NOR2_X1   g792(.A1(new_n189), .A2(G952), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n961), .A2(new_n966), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(G210), .A3(G902), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT56), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n521), .A2(new_n523), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(new_n526), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT55), .Z(new_n987));
  OAI21_X1  g801(.A(new_n980), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n984), .A2(new_n987), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n984), .A2(KEYINPUT120), .A3(new_n987), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G51));
  NAND2_X1  g807(.A1(new_n967), .A2(KEYINPUT121), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT121), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n961), .A2(new_n966), .A3(new_n995), .A4(new_n962), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n981), .A2(KEYINPUT54), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n360), .B(KEYINPUT57), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n777), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n981), .A2(G902), .A3(new_n856), .A4(new_n857), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n979), .B1(new_n1002), .B2(new_n1003), .ZN(G54));
  NAND4_X1  g818(.A1(new_n981), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n251), .A2(new_n259), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n1005), .A2(KEYINPUT122), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT122), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n979), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(G60));
  XNOR2_X1  g825(.A(new_n709), .B(KEYINPUT59), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n960), .B2(new_n967), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n705), .A2(new_n706), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n980), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1014), .A2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n998), .B2(new_n1017), .ZN(G63));
  INV_X1    g832(.A(KEYINPUT61), .ZN(new_n1019));
  INV_X1    g833(.A(new_n981), .ZN(new_n1020));
  XNOR2_X1  g834(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G217), .A2(G902), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n655), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n980), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n726), .A2(new_n728), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1020), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1019), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1027), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1029), .A2(KEYINPUT61), .A3(new_n980), .A4(new_n1024), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(G66));
  OAI21_X1  g845(.A(G953), .B1(new_n352), .B2(new_n506), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n805), .A2(new_n794), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1034), .A2(new_n678), .A3(new_n922), .A4(new_n931), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(new_n189), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n985), .B1(G898), .B2(new_n189), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1036), .B(new_n1037), .Z(G69));
  OAI22_X1  g852(.A1(new_n566), .A2(new_n567), .B1(KEYINPUT30), .B2(new_n571), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n222), .B1(new_n224), .B2(new_n221), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G900), .A2(G953), .ZN(new_n1042));
  AND3_X1   g856(.A1(new_n942), .A2(new_n743), .A3(new_n770), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1043), .A2(new_n843), .A3(new_n846), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n838), .A2(new_n943), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n866), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n874), .A2(new_n1046), .A3(new_n882), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1041), .B(new_n1042), .C1(new_n1047), .C2(G953), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n285), .A2(new_n712), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n839), .B1(new_n1049), .B2(new_n925), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n748), .B(new_n1050), .C1(new_n677), .C2(new_n675), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1051), .B(KEYINPUT125), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1043), .A2(new_n767), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1054));
  AND4_X1   g868(.A1(new_n874), .A2(new_n882), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1056), .B(KEYINPUT124), .ZN(new_n1057));
  AOI21_X1  g871(.A(G953), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1048), .B1(new_n1058), .B2(new_n1041), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1060));
  XOR2_X1   g874(.A(new_n1060), .B(KEYINPUT127), .Z(new_n1061));
  INV_X1    g875(.A(KEYINPUT126), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1061), .B1(new_n1048), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g878(.A(new_n1048), .B1(new_n1062), .B2(new_n1061), .C1(new_n1058), .C2(new_n1041), .ZN(new_n1065));
  AND2_X1   g879(.A1(new_n1064), .A2(new_n1065), .ZN(G72));
  NAND3_X1  g880(.A1(new_n1055), .A2(new_n754), .A3(new_n1057), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n753), .A2(new_n593), .ZN(new_n1068));
  OR2_X1    g882(.A1(new_n1047), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1035), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g884(.A(new_n754), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1071), .A2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g886(.A1(G472), .A2(G902), .ZN(new_n1073));
  XNOR2_X1  g887(.A(new_n1073), .B(KEYINPUT63), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n956), .A2(new_n959), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n979), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1070), .A2(new_n1078), .ZN(G57));
endmodule


