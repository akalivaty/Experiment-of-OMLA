//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1161, new_n1162, new_n1163, new_n1164, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n207), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n214), .B(new_n215), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(KEYINPUT1), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n244), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n248));
  AND2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n208), .B1(new_n203), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n209), .A2(G1), .ZN(new_n253));
  OR3_X1    g0053(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT70), .B1(new_n253), .B2(new_n217), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G150), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n250), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G50), .A2(G58), .ZN(new_n263));
  INV_X1    g0063(.A(G68), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n209), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n251), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n247), .A2(new_n248), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n256), .B(new_n266), .C1(G50), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT73), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(G1), .B(G13), .C1(new_n250), .C2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(G1698), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT67), .B(G223), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n276), .B1(new_n277), .B2(new_n274), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(new_n281), .B2(new_n280), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT66), .B(G41), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n244), .B(G274), .C1(new_n285), .C2(G45), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n273), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n283), .B(new_n286), .C1(new_n218), .C2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n269), .B(new_n270), .C1(new_n271), .C2(new_n289), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT72), .B(G200), .Z(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n268), .C1(G179), .C2(new_n289), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n259), .A2(new_n253), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT77), .Z(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(new_n252), .B1(new_n249), .B2(new_n259), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n251), .ZN(new_n304));
  INV_X1    g0104(.A(G58), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n264), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G58), .A2(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(G20), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT76), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(G159), .B2(new_n257), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT7), .B1(new_n313), .B2(new_n209), .ZN(new_n314));
  OR2_X1    g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  AND4_X1   g0116(.A1(KEYINPUT7), .A2(new_n315), .A3(new_n209), .A4(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n310), .B1(new_n264), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n304), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n310), .B(KEYINPUT16), .C1(new_n264), .C2(new_n318), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n303), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n286), .B1(new_n229), .B2(new_n288), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n218), .A2(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n274), .B(new_n326), .C1(G223), .C2(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G87), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n273), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n296), .B1(new_n325), .B2(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT78), .Z(new_n335));
  INV_X1    g0135(.A(KEYINPUT18), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n324), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n324), .B2(new_n335), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G190), .B2(new_n330), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n323), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n323), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G238), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n286), .B1(new_n349), .B2(new_n288), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n229), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n274), .B(new_n351), .C1(G226), .C2(G1698), .ZN(new_n352));
  AND3_X1   g0152(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n273), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G169), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n331), .C2(new_n359), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n267), .A2(G68), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n264), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n261), .B2(new_n277), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n251), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT11), .Z(new_n369));
  NOR2_X1   g0169(.A1(new_n253), .A2(new_n264), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n365), .B(new_n369), .C1(new_n252), .C2(new_n370), .ZN(new_n371));
  XOR2_X1   g0171(.A(new_n371), .B(KEYINPUT75), .Z(new_n372));
  NAND2_X1  g0172(.A1(new_n363), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n359), .A2(G200), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n371), .B(new_n374), .C1(new_n271), .C2(new_n359), .ZN(new_n375));
  INV_X1    g0175(.A(new_n259), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT71), .B1(new_n379), .B2(new_n260), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n251), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n253), .A2(new_n277), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n252), .A2(new_n384), .B1(new_n277), .B2(new_n249), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G232), .A2(G1698), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n275), .A2(G238), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n274), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n273), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(G107), .C2(new_n274), .ZN(new_n392));
  INV_X1    g0192(.A(G244), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n286), .C1(new_n393), .C2(new_n288), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n292), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n387), .B(new_n395), .C1(new_n271), .C2(new_n394), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(G179), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n296), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n386), .ZN(new_n399));
  AND4_X1   g0199(.A1(new_n373), .A2(new_n375), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  AND4_X1   g0200(.A1(new_n299), .A2(new_n339), .A3(new_n348), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n244), .A2(G33), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n267), .A2(new_n304), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G116), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n267), .A2(new_n219), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G283), .ZN(new_n407));
  INV_X1    g0207(.A(G97), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n209), .C1(G33), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT85), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n250), .A2(G97), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(KEYINPUT85), .A3(new_n209), .A4(new_n407), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n219), .A2(G20), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n251), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT84), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n411), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n251), .A2(KEYINPUT84), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n411), .A2(new_n413), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n416), .ZN(new_n421));
  AND4_X1   g0221(.A1(KEYINPUT20), .A2(new_n420), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n406), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n273), .A2(G274), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT5), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT66), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G41), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n244), .A2(G45), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(G41), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT5), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n438), .A2(KEYINPUT81), .A3(new_n433), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n426), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n274), .A2(G257), .A3(new_n275), .ZN(new_n442));
  INV_X1    g0242(.A(G303), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n274), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n391), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n434), .B(new_n424), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n273), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n440), .B(new_n445), .C1(new_n220), .C2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n423), .A2(new_n448), .A3(KEYINPUT21), .A4(G169), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT86), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n447), .A2(new_n220), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n432), .A2(new_n427), .A3(new_n434), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT81), .B1(new_n438), .B2(new_n433), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n425), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n296), .B1(new_n456), .B2(new_n445), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n423), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n423), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT21), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n448), .A2(new_n331), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n423), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(G190), .A3(new_n445), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n423), .B1(G200), .B2(new_n448), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n407), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  OAI211_X1 g0270(.A(G244), .B(new_n275), .C1(new_n311), .C2(new_n312), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n470), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n391), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n446), .A2(G257), .A3(new_n273), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n455), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n446), .A2(G257), .A3(new_n273), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT82), .B1(new_n440), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n249), .A2(new_n408), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n403), .B2(new_n408), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(G97), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT6), .A2(G97), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G107), .ZN(new_n491));
  AND2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NOR2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n488), .B(new_n491), .C1(new_n494), .C2(KEYINPUT6), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n314), .B2(new_n317), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n486), .B1(new_n498), .B2(new_n251), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n476), .A2(new_n469), .A3(new_n473), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n440), .B(new_n481), .C1(new_n500), .C2(new_n273), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT83), .B1(new_n501), .B2(new_n271), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n455), .A2(new_n478), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n477), .A2(new_n503), .A3(G190), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n484), .A2(new_n499), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n499), .B1(new_n501), .B2(new_n296), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n331), .B(new_n477), .C1(new_n480), .C2(new_n482), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n403), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n267), .B2(G107), .ZN(new_n514));
  AOI22_X1  g0314(.A1(G107), .A2(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n209), .B(G87), .C1(new_n311), .C2(new_n312), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT22), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT22), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n274), .A2(new_n519), .A3(new_n209), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n209), .B2(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n487), .A2(KEYINPUT23), .A3(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n260), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n521), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n516), .B1(new_n533), .B2(new_n251), .ZN(new_n534));
  AOI211_X1 g0334(.A(KEYINPUT24), .B(new_n527), .C1(new_n518), .C2(new_n520), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n521), .B2(new_n528), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n516), .B(new_n251), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n515), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n540));
  OAI211_X1 g0340(.A(G250), .B(new_n275), .C1(new_n311), .C2(new_n312), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n391), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n446), .A2(G264), .A3(new_n273), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR4_X1   g0346(.A1(new_n546), .A2(new_n455), .A3(KEYINPUT88), .A4(new_n331), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT88), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n546), .A2(new_n455), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G179), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n440), .A2(new_n545), .A3(new_n544), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G169), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n547), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n340), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n551), .B2(G190), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n515), .C1(new_n534), .C2(new_n538), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n511), .A2(new_n379), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT19), .B1(new_n353), .B2(new_n354), .ZN(new_n559));
  INV_X1    g0359(.A(G87), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n209), .B1(new_n560), .B2(new_n493), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n274), .A2(new_n209), .A3(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n260), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n251), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n249), .A2(new_n378), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n558), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G238), .B(new_n275), .C1(new_n311), .C2(new_n312), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n391), .ZN(new_n574));
  INV_X1    g0374(.A(G250), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n433), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G274), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n244), .A2(new_n577), .A3(G45), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n273), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n569), .B1(G179), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n573), .B2(new_n391), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(G169), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n581), .A2(G190), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(new_n292), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n267), .A2(new_n304), .A3(G87), .A4(new_n402), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n567), .A2(new_n568), .A3(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n582), .A2(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n554), .A2(new_n557), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n401), .A2(new_n467), .A3(new_n510), .A4(new_n593), .ZN(G372));
  NAND2_X1  g0394(.A1(new_n324), .A2(new_n335), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT18), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n324), .A2(new_n335), .A3(new_n336), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n399), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n375), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n373), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n348), .ZN(new_n602));
  INV_X1    g0402(.A(new_n295), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n298), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT91), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n507), .A2(new_n508), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n589), .A2(KEYINPUT90), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n567), .A2(new_n609), .A3(new_n568), .A4(new_n588), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n587), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n583), .A2(new_n331), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n569), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT89), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n581), .B2(new_n296), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n583), .A2(KEYINPUT89), .A3(G169), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n607), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT26), .B1(new_n509), .B2(new_n590), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n614), .A2(new_n618), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n554), .A2(new_n459), .A3(new_n463), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n506), .A2(new_n509), .A3(new_n557), .A4(new_n619), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n401), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT92), .ZN(G369));
  NAND3_X1  g0430(.A1(new_n244), .A2(new_n209), .A3(G13), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G343), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n423), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g0437(.A(new_n464), .B(new_n467), .S(new_n637), .Z(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n554), .A2(new_n557), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n539), .A2(new_n636), .ZN(new_n643));
  INV_X1    g0443(.A(new_n636), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n642), .A2(new_n643), .B1(new_n554), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n464), .A2(new_n644), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n554), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n644), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(G399));
  NAND2_X1  g0451(.A1(new_n284), .A2(new_n204), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n493), .A2(new_n560), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G116), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n654), .A3(G1), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n211), .B2(new_n652), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT28), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n607), .A2(new_n619), .A3(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n620), .B1(new_n509), .B2(new_n590), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n624), .B(new_n660), .C1(new_n625), .C2(new_n626), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n661), .A2(KEYINPUT93), .A3(new_n644), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT93), .B1(new_n661), .B2(new_n644), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT29), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n627), .A2(new_n644), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT29), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n546), .A2(new_n581), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n462), .A2(new_n477), .A3(new_n504), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n549), .A2(G179), .A3(new_n583), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n483), .A2(new_n672), .A3(new_n448), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n636), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT31), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n467), .A2(new_n510), .A3(new_n593), .A4(new_n644), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n664), .A2(new_n667), .B1(G330), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n657), .B1(new_n680), .B2(G1), .ZN(G364));
  NAND2_X1  g0481(.A1(new_n209), .A2(G13), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT94), .Z(new_n683));
  AOI21_X1  g0483(.A(new_n244), .B1(new_n683), .B2(G45), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n652), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n640), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(G330), .B2(new_n638), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n274), .A2(new_n204), .ZN(new_n690));
  INV_X1    g0490(.A(G355), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n690), .A2(new_n691), .B1(G116), .B2(new_n204), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n239), .A2(G45), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n313), .A2(new_n204), .ZN(new_n694));
  INV_X1    g0494(.A(G45), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n212), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(G20), .B1(KEYINPUT95), .B2(G169), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(KEYINPUT95), .A2(G169), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n208), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(G13), .A2(G33), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G20), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n687), .B1(new_n697), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n209), .A2(G190), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G179), .A2(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(G329), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n209), .A2(new_n331), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(G190), .A3(new_n340), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n274), .B(new_n712), .C1(G322), .C2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n291), .A2(new_n209), .A3(G179), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G303), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G283), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n271), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT97), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n713), .A2(G200), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(new_n726), .B2(new_n271), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n725), .A2(KEYINPUT97), .A3(G190), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT33), .B(G317), .Z(new_n730));
  OAI221_X1 g0530(.A(new_n721), .B1(new_n722), .B2(new_n723), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n708), .A2(G179), .A3(new_n340), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n209), .B1(new_n709), .B2(G190), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n725), .A2(new_n271), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(G326), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT98), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT96), .B(G159), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n711), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT32), .Z(new_n742));
  INV_X1    g0542(.A(new_n734), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n737), .A2(G50), .B1(G97), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n742), .B(new_n744), .C1(new_n264), .C2(new_n729), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n274), .B1(new_n732), .B2(new_n277), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(G58), .B2(new_n715), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n747), .B1(new_n723), .B2(new_n487), .C1(new_n560), .C2(new_n718), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n731), .A2(new_n739), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n707), .B1(new_n749), .B2(new_n701), .ZN(new_n750));
  INV_X1    g0550(.A(new_n704), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n638), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n689), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(G396));
  NAND2_X1  g0554(.A1(new_n386), .A2(new_n636), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n599), .B1(new_n396), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n399), .A2(new_n636), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n665), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n627), .A2(new_n644), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n679), .A2(G330), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n687), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n701), .A2(new_n702), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n686), .B(new_n685), .C1(new_n277), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n701), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n560), .A2(new_n723), .B1(new_n718), .B2(new_n487), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n729), .A2(new_n722), .ZN(new_n770));
  INV_X1    g0570(.A(new_n732), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G116), .B1(new_n711), .B2(G311), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n313), .C1(new_n735), .C2(new_n714), .ZN(new_n773));
  INV_X1    g0573(.A(new_n737), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n774), .A2(new_n443), .B1(new_n734), .B2(new_n408), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n769), .A2(new_n770), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n313), .B1(new_n711), .B2(G132), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n217), .A2(new_n718), .B1(new_n723), .B2(new_n264), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n777), .B1(new_n305), .B2(new_n734), .C1(new_n778), .C2(KEYINPUT99), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(KEYINPUT99), .B2(new_n778), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G143), .A2(new_n715), .B1(new_n771), .B2(new_n740), .ZN(new_n781));
  INV_X1    g0581(.A(G137), .ZN(new_n782));
  INV_X1    g0582(.A(G150), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n774), .C1(new_n729), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT34), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n776), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n767), .B1(new_n768), .B2(new_n786), .C1(new_n758), .C2(new_n703), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n765), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G384));
  OR2_X1    g0589(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n790), .A2(G116), .A3(new_n210), .A4(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT36), .Z(new_n793));
  OAI211_X1 g0593(.A(new_n212), .B(G77), .C1(new_n305), .C2(new_n264), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n217), .A2(G68), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n244), .B(G13), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT38), .ZN(new_n798));
  INV_X1    g0598(.A(new_n634), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n324), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n339), .B2(new_n348), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n595), .A2(new_n800), .A3(new_n343), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT37), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n595), .A2(new_n800), .A3(KEYINPUT37), .A4(new_n343), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n800), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n598), .B2(new_n347), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n809), .A2(KEYINPUT38), .A3(new_n805), .A4(new_n804), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT39), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(KEYINPUT39), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n363), .A2(new_n372), .A3(new_n644), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT101), .Z(new_n817));
  OAI22_X1  g0617(.A1(new_n815), .A2(new_n817), .B1(new_n339), .B2(new_n799), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n807), .A2(new_n810), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n373), .A2(new_n375), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(new_n372), .A3(new_n636), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n372), .A2(new_n636), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n373), .A2(new_n822), .A3(new_n375), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n757), .B(KEYINPUT100), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n761), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n818), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n401), .A2(new_n667), .A3(new_n664), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n606), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n830), .B(new_n832), .Z(new_n833));
  INV_X1    g0633(.A(G330), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT102), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n679), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n759), .B1(new_n821), .B2(new_n823), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n811), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT40), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(KEYINPUT40), .A3(new_n811), .A4(new_n837), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n401), .A2(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n244), .B2(new_n683), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n833), .A2(new_n847), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n797), .B1(new_n849), .B2(new_n850), .ZN(G367));
  OAI21_X1  g0651(.A(new_n510), .B1(new_n499), .B2(new_n644), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT103), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n509), .B1(new_n853), .B2(new_n554), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n644), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n509), .B2(new_n644), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n648), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT42), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n859), .A2(new_n860), .B1(new_n858), .B2(new_n857), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n619), .B1(new_n611), .B2(new_n644), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n624), .A2(new_n611), .A3(new_n644), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n861), .A2(new_n862), .B1(KEYINPUT43), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT43), .B2(new_n865), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n856), .A2(new_n640), .A3(new_n645), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT43), .ZN(new_n869));
  INV_X1    g0669(.A(new_n865), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n861), .A2(new_n862), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n868), .B1(new_n867), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n652), .B(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT106), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(KEYINPUT44), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n856), .A2(new_n650), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT44), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(KEYINPUT106), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n878), .B(KEYINPUT44), .C1(new_n856), .C2(new_n650), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n650), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT45), .B1(new_n856), .B2(new_n650), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OR3_X1    g0687(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n646), .ZN(new_n888));
  INV_X1    g0688(.A(new_n648), .ZN(new_n889));
  INV_X1    g0689(.A(new_n647), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n645), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n639), .B(new_n891), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n680), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n646), .B1(new_n887), .B2(KEYINPUT107), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n877), .B1(new_n899), .B2(new_n680), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n874), .B1(new_n900), .B2(new_n685), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n235), .A2(new_n694), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n705), .B1(new_n204), .B2(new_n378), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n687), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT109), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n774), .A2(new_n733), .B1(new_n734), .B2(new_n487), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n313), .B1(new_n732), .B2(new_n722), .ZN(new_n907));
  INV_X1    g0707(.A(G317), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n714), .A2(new_n443), .B1(new_n710), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n910), .B1(new_n408), .B2(new_n723), .C1(new_n735), .C2(new_n729), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n718), .A2(new_n219), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT46), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n714), .A2(new_n783), .B1(new_n734), .B2(new_n264), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(G143), .B2(new_n737), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT110), .ZN(new_n916));
  INV_X1    g0716(.A(new_n729), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n740), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n719), .A2(G58), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n274), .B1(new_n710), .B2(new_n782), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(G50), .B2(new_n771), .ZN(new_n921));
  INV_X1    g0721(.A(new_n723), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G77), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n918), .A2(new_n919), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n911), .A2(new_n913), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT47), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n701), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n905), .B1(new_n865), .B2(new_n751), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n901), .A2(new_n930), .ZN(G387));
  OAI211_X1 g0731(.A(new_n896), .B(new_n686), .C1(new_n680), .C2(new_n892), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n645), .A2(new_n751), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n690), .A2(new_n654), .B1(G107), .B2(new_n204), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT111), .Z(new_n935));
  OR2_X1    g0735(.A1(new_n232), .A2(new_n695), .ZN(new_n936));
  INV_X1    g0736(.A(new_n654), .ZN(new_n937));
  AOI211_X1 g0737(.A(G45), .B(new_n937), .C1(G68), .C2(G77), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n259), .A2(G50), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n694), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n935), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n687), .B1(new_n942), .B2(new_n706), .ZN(new_n943));
  INV_X1    g0743(.A(G159), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n774), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT112), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n718), .A2(new_n277), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n922), .A2(G97), .B1(new_n945), .B2(KEYINPUT112), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n917), .A2(new_n376), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n714), .A2(new_n217), .B1(new_n732), .B2(new_n264), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n734), .A2(new_n378), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n274), .B1(new_n710), .B2(new_n783), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n274), .B1(new_n711), .B2(G326), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n718), .A2(new_n735), .B1(new_n722), .B2(new_n734), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G317), .A2(new_n715), .B1(new_n771), .B2(G303), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT113), .B(G322), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n958), .B1(new_n774), .B2(new_n959), .C1(new_n729), .C2(new_n733), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT48), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT49), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n956), .B1(new_n219), .B2(new_n723), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n955), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n943), .B1(new_n967), .B2(new_n701), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n892), .A2(new_n685), .B1(new_n933), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n932), .A2(new_n969), .ZN(G393));
  XNOR2_X1  g0770(.A(new_n886), .B(new_n646), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n899), .B(new_n686), .C1(new_n897), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n856), .A2(new_n751), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n242), .A2(new_n694), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n705), .B1(new_n408), .B2(new_n204), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n687), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT52), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n774), .A2(new_n908), .B1(new_n733), .B2(new_n714), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n917), .A2(G303), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G107), .A2(new_n922), .B1(new_n719), .B2(G283), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n710), .A2(new_n959), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n313), .B1(new_n732), .B2(new_n735), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(G116), .C2(new_n743), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n978), .A2(new_n977), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n980), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G68), .A2(new_n719), .B1(new_n922), .B2(G87), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n734), .A2(new_n277), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n274), .B1(new_n732), .B2(new_n259), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G143), .C2(new_n711), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n989), .C1(new_n217), .C2(new_n729), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G150), .A2(new_n737), .B1(new_n715), .B2(G159), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT51), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n985), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n976), .B1(new_n993), .B2(new_n701), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n971), .A2(new_n685), .B1(new_n973), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n972), .A2(new_n995), .ZN(G390));
  AOI21_X1  g0796(.A(new_n703), .B1(new_n813), .B2(new_n814), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n771), .A2(G97), .B1(new_n711), .B2(G294), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n313), .C1(new_n219), .C2(new_n714), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n987), .B(new_n999), .C1(G283), .C2(new_n737), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G68), .A2(new_n922), .B1(new_n719), .B2(G87), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n487), .C2(new_n729), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n719), .A2(G150), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT53), .ZN(new_n1004));
  INV_X1    g0804(.A(G132), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n274), .B1(new_n714), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(G128), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n774), .A2(new_n1007), .B1(new_n734), .B2(new_n944), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(G125), .C2(new_n711), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT54), .B(G143), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT118), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n922), .A2(G50), .B1(new_n771), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n782), .C2(new_n729), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1002), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n701), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n766), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n687), .C1(new_n376), .C2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n997), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n828), .A2(new_n817), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n815), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n824), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n679), .A2(G330), .A3(new_n758), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n661), .A2(new_n644), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT93), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n661), .A2(KEYINPUT93), .A3(new_n644), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n759), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT114), .B1(new_n1029), .B2(new_n825), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n758), .B1(new_n662), .B2(new_n663), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT114), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n826), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n824), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT115), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n811), .A2(new_n817), .ZN(new_n1036));
  AND3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1035), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1020), .B(new_n1024), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n815), .A2(new_n1019), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT115), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n842), .A2(G330), .A3(new_n837), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT117), .B1(new_n1046), .B2(new_n684), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1020), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1045), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT117), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n685), .A4(new_n1039), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1018), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT116), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n401), .A2(new_n842), .A3(G330), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n606), .A2(new_n1055), .A3(new_n831), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n827), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n836), .A2(G330), .A3(new_n758), .A4(new_n838), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n1021), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1024), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1056), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1046), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1039), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1066));
  AND4_X1   g0866(.A1(new_n1054), .A2(new_n1065), .A3(new_n686), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n652), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1054), .B1(new_n1068), .B2(new_n1066), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1053), .B1(new_n1067), .B2(new_n1069), .ZN(G378));
  XNOR2_X1  g0870(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n268), .A2(new_n799), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n299), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n299), .A2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1076), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n841), .A2(G330), .A3(new_n843), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(new_n843), .A3(G330), .A4(new_n841), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n830), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n830), .A3(new_n1084), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n685), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1081), .A2(new_n702), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n687), .B1(G50), .B2(new_n1016), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n723), .A2(new_n305), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT120), .Z(new_n1094));
  NAND2_X1  g0894(.A1(new_n917), .A2(G97), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n737), .A2(G116), .B1(G68), .B2(new_n743), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n313), .B(new_n284), .C1(new_n732), .C2(new_n378), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n714), .A2(new_n487), .B1(new_n710), .B2(new_n722), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n947), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1094), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT58), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n734), .A2(new_n783), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n714), .A2(new_n1007), .B1(new_n732), .B2(new_n782), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G125), .C2(new_n737), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n719), .A2(new_n1011), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n1005), .C2(new_n729), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n922), .A2(new_n740), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G33), .B(G41), .C1(new_n711), .C2(G124), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1101), .A2(KEYINPUT58), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n217), .B1(G33), .B2(G41), .C1(new_n285), .C2(new_n274), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT119), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1102), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1092), .B1(new_n1116), .B2(new_n701), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1091), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1090), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1056), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1066), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1089), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT57), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n652), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT121), .Z(G375));
  NAND3_X1  g0928(.A1(new_n1058), .A2(new_n1056), .A3(new_n1062), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1064), .A2(new_n876), .A3(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT122), .Z(new_n1131));
  AOI21_X1  g0931(.A(new_n684), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT123), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n687), .B1(G68), .B2(new_n1016), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n771), .A2(G107), .B1(new_n711), .B2(G303), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n313), .C1(new_n722), .C2(new_n714), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n952), .B(new_n1137), .C1(G294), .C2(new_n737), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G77), .A2(new_n922), .B1(new_n719), .B2(G97), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n219), .C2(new_n729), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n274), .B1(new_n710), .B2(new_n1007), .C1(new_n714), .C2(new_n782), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G132), .B2(new_n737), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1094), .B(new_n1142), .C1(new_n944), .C2(new_n718), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT124), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n732), .A2(new_n783), .B1(new_n734), .B2(new_n217), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n917), .A2(new_n1011), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1140), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1135), .B1(new_n1148), .B2(new_n701), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n824), .B2(new_n703), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1133), .A2(KEYINPUT123), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1134), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1131), .A2(new_n1152), .ZN(G381));
  NAND2_X1  g0953(.A1(new_n1068), .A2(new_n1066), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1053), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(G393), .A2(G396), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1131), .A2(new_n788), .A3(new_n1152), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G390), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n901), .A3(new_n930), .ZN(new_n1159));
  OR4_X1    g0959(.A1(G375), .A2(new_n1155), .A3(new_n1157), .A4(new_n1159), .ZN(G407));
  INV_X1    g0960(.A(new_n1155), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n635), .A2(G213), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G407), .B(G213), .C1(G375), .C2(new_n1164), .ZN(G409));
  NOR2_X1   g0965(.A1(new_n1122), .A2(new_n877), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1090), .A2(KEYINPUT126), .A3(new_n1118), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT126), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n684), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1118), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1161), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT125), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1127), .A2(G378), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1127), .B2(G378), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n686), .B(new_n1064), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1152), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n788), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1152), .A2(G384), .A3(new_n1181), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1177), .A2(new_n1162), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT62), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT61), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1163), .A2(G2897), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1185), .B(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1127), .A2(G378), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT125), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1127), .A2(G378), .A3(new_n1174), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1172), .A2(new_n1166), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1193), .A2(new_n1194), .B1(new_n1161), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1196), .B2(new_n1163), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT62), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1177), .A2(new_n1198), .A3(new_n1162), .A4(new_n1186), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1188), .A2(new_n1189), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n753), .B1(new_n932), .B2(new_n969), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1156), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1159), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1158), .B1(new_n901), .B2(new_n930), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(G387), .A2(G390), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1202), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1159), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1200), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT63), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1187), .B2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1177), .A2(KEYINPUT63), .A3(new_n1162), .A4(new_n1186), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1212), .A2(new_n1189), .A3(new_n1213), .A4(new_n1197), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(G405));
  AND2_X1   g1015(.A1(G375), .A2(new_n1161), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1216), .A2(new_n1217), .B1(KEYINPUT127), .B2(new_n1186), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1205), .A2(new_n1208), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1218), .B(new_n1222), .ZN(G402));
endmodule


