//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G116), .B(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT69), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n199));
  OAI21_X1  g013(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n204), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n205), .B2(new_n210), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n193), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n213), .B1(new_n209), .B2(new_n212), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n195), .A2(new_n197), .A3(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n218), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n222), .B(new_n224), .C1(new_n225), .C2(new_n220), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(new_n226), .A3(new_n228), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(KEYINPUT81), .A3(new_n231), .A4(KEYINPUT6), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT66), .B1(new_n237), .B2(G143), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT64), .A2(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT64), .A2(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n241), .B2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NOR4_X1   g057(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT66), .A4(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n236), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n243), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT65), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT64), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT64), .A2(G146), .ZN(new_n255));
  AOI21_X1  g069(.A(G143), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n250), .C1(new_n256), .C2(new_n246), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n245), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(G143), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n248), .B1(G128), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n238), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n241), .A2(new_n268), .A3(G143), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G125), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n263), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n259), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G224), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT83), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n259), .B2(new_n273), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n281), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n279), .B1(new_n284), .B2(new_n275), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n235), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT84), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n259), .A2(new_n288), .B1(KEYINPUT7), .B2(new_n279), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n259), .A2(new_n273), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n214), .A2(new_n215), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n202), .A2(new_n218), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n228), .B(KEYINPUT8), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n196), .A2(KEYINPUT5), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n218), .B1(new_n296), .B2(new_n200), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n216), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n291), .A2(new_n231), .A3(new_n292), .A4(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n188), .B1(new_n287), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n292), .A2(new_n231), .A3(new_n299), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n305), .B2(new_n291), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n234), .B(new_n232), .C1(new_n285), .C2(new_n282), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n187), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT85), .A4(new_n187), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G128), .B1(new_n246), .B2(new_n264), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n267), .A2(new_n269), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n293), .B1(new_n271), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n222), .B1(new_n225), .B2(new_n220), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(new_n258), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n330), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n263), .A2(new_n271), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n323), .A2(new_n325), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G140), .ZN(new_n341));
  INV_X1    g155(.A(G227), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G953), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT80), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(KEYINPUT80), .A3(new_n345), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n338), .A2(new_n216), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n336), .B1(new_n349), .B2(new_n320), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n323), .A2(new_n325), .A3(new_n339), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n336), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n340), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n347), .A2(new_n354), .B1(new_n357), .B2(new_n345), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n301), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n301), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n340), .B1(new_n353), .B2(new_n352), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(new_n344), .B1(new_n356), .B2(new_n346), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(G469), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n317), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G237), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n277), .A3(G214), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(KEYINPUT86), .B2(new_n243), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT86), .B(G143), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n370), .B2(G131), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n373), .A3(G131), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n272), .A3(G140), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT16), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n272), .B2(G140), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n237), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n378), .A2(KEYINPUT19), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n381), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(KEYINPUT19), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n247), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n370), .A2(G131), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n371), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n241), .A2(new_n378), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n388), .B2(new_n237), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n393), .B2(new_n370), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n377), .A2(new_n390), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  INV_X1    g220(.A(new_n376), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n406), .B(new_n371), .C1(new_n407), .C2(new_n374), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n382), .A2(new_n237), .A3(new_n384), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n385), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n386), .A2(KEYINPUT89), .A3(new_n410), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n376), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n396), .A2(new_n399), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n403), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT20), .B1(new_n405), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT90), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  INV_X1    g236(.A(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n405), .B2(new_n417), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n415), .A2(new_n416), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n404), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n301), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G475), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G234), .A2(G237), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(G952), .A3(new_n277), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(G902), .A3(G953), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n434), .B(KEYINPUT92), .Z(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(G107), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT91), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n203), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G128), .B(G143), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n445));
  INV_X1    g259(.A(G128), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n446), .A2(KEYINPUT13), .A3(G143), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n327), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n445), .A2(new_n448), .B1(new_n327), .B2(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n444), .B(new_n327), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n438), .ZN(new_n453));
  OAI211_X1 g267(.A(G107), .B(new_n452), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(new_n454), .C1(G107), .C2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n315), .A2(new_n457), .A3(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n455), .A3(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n301), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n431), .A2(new_n437), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n314), .A2(new_n365), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G472), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT67), .B1(new_n329), .B2(G134), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n327), .A3(G137), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n329), .A2(G134), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G131), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n477), .A2(new_n335), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n262), .B2(new_n270), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n245), .A2(new_n252), .A3(new_n336), .A4(new_n257), .ZN(new_n480));
  INV_X1    g294(.A(new_n224), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n483), .A2(KEYINPUT28), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(KEYINPUT73), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n224), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n479), .A2(new_n480), .A3(new_n488), .A4(new_n481), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n495));
  INV_X1    g309(.A(G210), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(G237), .A3(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n493), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n483), .A2(KEYINPUT28), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(new_n504), .A3(new_n487), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(new_n501), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT30), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n479), .A2(new_n480), .A3(new_n509), .A4(KEYINPUT30), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n479), .C2(new_n480), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n486), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n511), .B(new_n224), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n516), .A2(new_n482), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n506), .B(new_n494), .C1(new_n517), .C2(new_n500), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n471), .B1(new_n503), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n500), .A3(new_n482), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT31), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n516), .A2(new_n524), .A3(new_n500), .A4(new_n482), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n505), .A2(new_n501), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n471), .A3(new_n301), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n519), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n529), .A2(KEYINPUT32), .A3(new_n471), .A4(new_n301), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT72), .B1(new_n520), .B2(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n526), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n471), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT77), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n189), .B2(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n446), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(new_n546), .C1(G119), .C2(new_n446), .ZN(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT24), .B(G110), .Z(new_n549));
  AOI22_X1  g363(.A1(new_n547), .A2(G110), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n411), .B2(new_n385), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n547), .A2(G110), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n386), .A2(new_n397), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT76), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT22), .B(G137), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n551), .B2(new_n553), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n543), .B1(new_n560), .B2(G902), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT25), .B(new_n301), .C1(new_n558), .C2(new_n559), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n457), .B1(G234), .B2(new_n301), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(G902), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n558), .B2(new_n559), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n541), .A2(new_n542), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n542), .B1(new_n541), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n470), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  AOI21_X1  g388(.A(new_n471), .B1(new_n529), .B2(new_n301), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n530), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n365), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n569), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n463), .A2(new_n464), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT93), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n463), .A2(KEYINPUT93), .A3(new_n464), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n462), .B(KEYINPUT33), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n464), .A2(G902), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n425), .B2(new_n430), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n303), .A2(new_n308), .ZN(new_n590));
  INV_X1    g404(.A(new_n437), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n312), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n581), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT34), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n312), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n430), .A2(new_n468), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT94), .B1(new_n424), .B2(new_n422), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n418), .A2(new_n419), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n424), .A2(KEYINPUT94), .A3(new_n422), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT95), .A3(new_n599), .A4(new_n600), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n597), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n581), .A2(new_n437), .A3(new_n596), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT35), .B(G107), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NAND2_X1  g424(.A1(new_n551), .A2(new_n553), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(new_n567), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n565), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n470), .A2(new_n578), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G12));
  INV_X1    g433(.A(new_n596), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n435), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(KEYINPUT96), .ZN(new_n623));
  INV_X1    g437(.A(new_n433), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n622), .B2(KEYINPUT96), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AND4_X1   g441(.A1(new_n620), .A2(new_n606), .A3(new_n616), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n541), .A2(new_n628), .A3(new_n365), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G128), .ZN(G30));
  XOR2_X1   g444(.A(new_n626), .B(KEYINPUT39), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n365), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n311), .B(KEYINPUT38), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n425), .A2(new_n430), .B1(new_n467), .B2(new_n466), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n615), .A3(new_n312), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n535), .A2(new_n540), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n517), .A2(new_n501), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n491), .B2(new_n501), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n471), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n530), .B2(new_n531), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n637), .B(new_n644), .C1(KEYINPUT40), .C2(new_n632), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G143), .ZN(G45));
  AOI211_X1 g460(.A(new_n626), .B(new_n588), .C1(new_n430), .C2(new_n425), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n648), .A2(new_n596), .A3(new_n615), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n541), .A2(new_n365), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT97), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n541), .A2(new_n649), .A3(new_n652), .A4(new_n365), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G146), .ZN(G48));
  NAND2_X1  g469(.A1(new_n358), .A2(new_n301), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G469), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n316), .A3(new_n360), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n592), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n541), .A2(new_n570), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n596), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n541), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n606), .A2(new_n570), .A3(new_n591), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G116), .ZN(G18));
  AND2_X1   g482(.A1(new_n469), .A2(new_n616), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G119), .ZN(G21));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n493), .A2(new_n501), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n521), .A2(new_n525), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(G472), .A2(G902), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n674), .A2(new_n672), .A3(new_n675), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n575), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n635), .A2(new_n312), .A3(new_n590), .A4(new_n591), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n658), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n680), .A3(new_n570), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G122), .ZN(G24));
  NOR4_X1   g496(.A1(new_n575), .A2(new_n677), .A3(new_n615), .A4(new_n676), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n647), .A3(new_n663), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n313), .B1(new_n309), .B2(new_n310), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n365), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n541), .A2(new_n570), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n686), .B1(new_n690), .B2(new_n648), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n688), .A2(new_n686), .A3(new_n648), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n569), .B1(new_n532), .B2(new_n533), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT99), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT99), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n691), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G131), .ZN(G33));
  NOR2_X1   g512(.A1(new_n607), .A2(new_n626), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n541), .A2(new_n699), .A3(new_n570), .A4(new_n689), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G134), .ZN(G36));
  INV_X1    g515(.A(new_n360), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n363), .A2(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n363), .A2(KEYINPUT45), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT100), .B1(new_n363), .B2(KEYINPUT45), .ZN(new_n707));
  OAI211_X1 g521(.A(G469), .B(new_n703), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n361), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(KEYINPUT46), .A3(new_n709), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n317), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n687), .B(KEYINPUT101), .Z(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n631), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n588), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n430), .A3(new_n425), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT43), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n615), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(KEYINPUT44), .A3(new_n577), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT44), .B1(new_n720), .B2(new_n577), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n716), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n329), .ZN(G39));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n714), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n728), .B1(new_n714), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n687), .A2(new_n569), .A3(new_n647), .ZN(new_n732));
  OR3_X1    g546(.A1(new_n541), .A2(KEYINPUT103), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT103), .B1(new_n541), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G140), .ZN(G42));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n629), .A2(new_n684), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n653), .B2(new_n651), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n620), .A2(new_n635), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n615), .A2(new_n627), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n579), .A2(KEYINPUT107), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT107), .B1(new_n579), .B2(new_n742), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n644), .A2(new_n741), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n629), .A2(new_n684), .ZN(new_n747));
  AND4_X1   g561(.A1(KEYINPUT52), .A2(new_n654), .A3(new_n747), .A4(new_n745), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n541), .B(new_n663), .C1(new_n666), .C2(new_n669), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n660), .A3(new_n681), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n660), .A4(new_n681), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n700), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT99), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n694), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n758), .B2(new_n691), .ZN(new_n759));
  INV_X1    g573(.A(new_n589), .ZN(new_n760));
  INV_X1    g574(.A(new_n425), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n597), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n591), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n578), .A2(new_n763), .A3(new_n314), .A4(new_n580), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n617), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n541), .A2(new_n570), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT77), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n541), .A2(new_n542), .A3(new_n570), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n769), .B2(new_n470), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n603), .A2(new_n605), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n468), .A2(new_n626), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n430), .B(new_n772), .C1(new_n565), .C2(new_n614), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n365), .A2(new_n687), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n687), .A2(new_n365), .A3(new_n647), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n541), .A2(new_n775), .B1(new_n683), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n755), .A2(new_n759), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n738), .B1(new_n749), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n777), .A2(new_n700), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n764), .A2(new_n617), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n573), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n573), .A2(new_n781), .A3(new_n782), .A4(KEYINPUT108), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n654), .A2(new_n745), .A3(new_n747), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n740), .A2(KEYINPUT52), .A3(new_n745), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n660), .A2(new_n681), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n750), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n796));
  AND4_X1   g610(.A1(KEYINPUT53), .A2(new_n795), .A3(new_n697), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n787), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n779), .A2(new_n780), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT106), .B1(new_n793), .B2(new_n750), .ZN(new_n800));
  INV_X1    g614(.A(new_n754), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n770), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n697), .A2(new_n700), .A3(new_n777), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n780), .B1(new_n779), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT110), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n749), .A2(new_n778), .A3(new_n738), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT53), .B1(new_n804), .B2(new_n792), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n779), .A2(new_n780), .A3(new_n798), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n658), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n687), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT116), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n816), .A2(new_n569), .A3(new_n624), .A4(new_n644), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n589), .ZN(new_n818));
  INV_X1    g632(.A(G952), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n678), .A2(new_n570), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n719), .A2(new_n624), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n819), .B(G953), .C1(new_n823), .C2(new_n663), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n816), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n693), .A3(new_n821), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT48), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n827), .B2(new_n830), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n825), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n431), .A2(new_n717), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n817), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n817), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n826), .A2(new_n683), .A3(new_n821), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n657), .A2(new_n360), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n316), .B1(new_n842), .B2(KEYINPUT112), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(KEYINPUT112), .B2(new_n842), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n730), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n823), .A2(new_n715), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n634), .A2(new_n313), .A3(new_n814), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n822), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT50), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(KEYINPUT51), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n834), .B1(new_n841), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n844), .B(KEYINPUT113), .Z(new_n855));
  OAI21_X1  g669(.A(new_n846), .B1(new_n731), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n851), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n854), .B(new_n856), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n807), .A2(new_n813), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n819), .A2(new_n277), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n644), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n842), .A2(KEYINPUT49), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT104), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n570), .A2(new_n316), .A3(new_n312), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n718), .B(new_n869), .C1(KEYINPUT49), .C2(new_n842), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n866), .A2(new_n634), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n865), .A2(new_n872), .ZN(G75));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n779), .A2(new_n798), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(G902), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT119), .B(new_n874), .C1(new_n876), .C2(new_n496), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n277), .A2(G952), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT120), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n286), .A2(new_n235), .A3(new_n283), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n307), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n301), .B1(new_n779), .B2(new_n798), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n886), .B2(KEYINPUT119), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n874), .B1(new_n876), .B2(new_n496), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n883), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n880), .B1(new_n887), .B2(new_n890), .ZN(G51));
  XNOR2_X1  g705(.A(new_n358), .B(KEYINPUT121), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n780), .B1(new_n779), .B2(new_n798), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n799), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n361), .B(KEYINPUT57), .Z(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n876), .A2(new_n708), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n878), .B1(new_n896), .B2(new_n897), .ZN(G54));
  NAND3_X1  g712(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n405), .A2(new_n417), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n878), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n586), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n879), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n799), .A2(new_n806), .A3(KEYINPUT110), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n811), .B1(new_n810), .B2(new_n812), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n586), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(G63));
  INV_X1    g728(.A(new_n879), .ZN(new_n915));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  AND3_X1   g731(.A1(new_n787), .A2(new_n792), .A3(new_n797), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n809), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n919), .B2(new_n560), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n613), .B(KEYINPUT123), .Z(new_n921));
  OAI211_X1 g735(.A(new_n917), .B(new_n921), .C1(new_n809), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n875), .A2(new_n924), .A3(new_n917), .A4(new_n921), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n920), .A2(KEYINPUT61), .A3(new_n922), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  INV_X1    g744(.A(G224), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n436), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n802), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n235), .B1(G898), .B2(new_n277), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  AOI21_X1  g750(.A(new_n730), .B1(new_n734), .B2(new_n733), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n723), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n740), .B(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n714), .A2(new_n631), .A3(new_n741), .A4(new_n693), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n938), .A2(new_n759), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n277), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n515), .A2(new_n512), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n508), .B2(new_n510), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n389), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n342), .B2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n621), .B1(new_n946), .B2(new_n342), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n940), .A2(new_n645), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n940), .A2(new_n645), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n762), .A2(new_n687), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n632), .B(new_n956), .C1(new_n767), .C2(new_n768), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n937), .A2(new_n723), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n953), .A2(new_n961), .A3(new_n955), .A4(new_n958), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n946), .A2(new_n277), .ZN(new_n964));
  OAI221_X1 g778(.A(new_n948), .B1(new_n277), .B2(new_n949), .C1(new_n963), .C2(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n942), .B2(new_n802), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n517), .A2(new_n501), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n878), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n520), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n517), .A2(new_n500), .ZN(new_n972));
  OAI221_X1 g786(.A(new_n967), .B1(new_n971), .B2(new_n972), .C1(new_n808), .C2(new_n809), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n960), .A2(new_n933), .A3(new_n962), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n976), .B2(new_n639), .ZN(G57));
endmodule


