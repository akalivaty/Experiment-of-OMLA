//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT65), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT67), .B(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n209), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  INV_X1    g0026(.A(new_n202), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n214), .B1(KEYINPUT1), .B2(new_n223), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n224), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n204), .A2(new_n209), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n209), .A2(new_n249), .A3(KEYINPUT70), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT70), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G20), .B2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n209), .A2(G33), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n247), .B1(new_n248), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n208), .A2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT71), .Z(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n263), .A2(new_n209), .A3(G1), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n247), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n262), .A2(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n259), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT72), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT68), .B1(new_n273), .B2(new_n224), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G1), .A4(G13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n272), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n274), .A2(new_n277), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(new_n270), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n281), .B2(G226), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(G1698), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT69), .B(G223), .Z(new_n287));
  OAI221_X1 g0087(.A(new_n285), .B1(new_n205), .B2(new_n283), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n273), .A2(new_n224), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n259), .A2(new_n267), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n294), .B2(KEYINPUT73), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n269), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n269), .B2(new_n297), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n291), .A2(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n296), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n291), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n300), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n254), .A2(new_n266), .ZN(new_n307));
  INV_X1    g0107(.A(new_n215), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n308), .A2(new_n209), .B1(new_n205), .B2(new_n257), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n247), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n265), .A2(G68), .A3(new_n260), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n263), .A2(G1), .ZN(new_n315));
  AND4_X1   g0115(.A1(KEYINPUT12), .A2(new_n215), .A3(G20), .A4(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G68), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT12), .B1(new_n264), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n283), .A2(G226), .A3(new_n284), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n289), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n274), .A2(G238), .A3(new_n277), .A4(new_n270), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n329), .B2(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n320), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT74), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT74), .A4(new_n331), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n334), .A2(G179), .A3(new_n332), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n336), .A2(new_n337), .A3(new_n343), .A4(G169), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n320), .B(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n265), .A2(G77), .A3(new_n260), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n315), .A2(G20), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n257), .B1(new_n209), .B2(new_n205), .ZN(new_n351));
  INV_X1    g0151(.A(new_n256), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n253), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n247), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n348), .B1(G77), .B2(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n279), .B1(new_n281), .B2(G244), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n358), .B2(new_n283), .C1(new_n286), .C2(new_n216), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n289), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(G200), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n321), .B2(new_n361), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n304), .A3(new_n360), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n355), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n306), .A2(new_n339), .A3(new_n347), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n283), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G33), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G68), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n227), .B1(new_n215), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n253), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n383), .A2(new_n247), .ZN(new_n384));
  INV_X1    g0184(.A(new_n378), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n382), .B1(new_n385), .B2(new_n215), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n265), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n352), .A2(new_n260), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n390), .A2(new_n391), .B1(new_n349), .B2(new_n352), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT78), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n270), .A2(G232), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n280), .B(new_n397), .C1(new_n272), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n274), .A3(new_n277), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n278), .A3(KEYINPUT76), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n373), .A2(new_n375), .A3(G226), .A4(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n373), .A2(new_n375), .A3(G223), .A4(new_n284), .ZN(new_n403));
  INV_X1    g0203(.A(G87), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n403), .C1(new_n249), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n289), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT77), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT77), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n399), .A2(new_n401), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n293), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n407), .A2(G190), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n396), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(G200), .B1(new_n408), .B2(new_n410), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n395), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n407), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n411), .A2(new_n364), .B1(new_n304), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n422), .A2(new_n394), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n422), .B2(new_n394), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n412), .A2(new_n396), .A3(new_n414), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT78), .B1(new_n416), .B2(new_n413), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n394), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT17), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n420), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n370), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n289), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n373), .A2(new_n375), .A3(G264), .A4(G1698), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n373), .A2(new_n375), .A3(G257), .A4(new_n284), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT83), .B(G303), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n434), .B(new_n435), .C1(new_n283), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT84), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT83), .B(G303), .Z(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n376), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT84), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n434), .A4(new_n435), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n433), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(new_n274), .A3(G270), .A4(new_n277), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n274), .A2(new_n451), .A3(new_n452), .A4(new_n277), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n209), .C1(G33), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n247), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n349), .A2(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n208), .A2(G33), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n354), .A2(new_n349), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G169), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT21), .B1(new_n455), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n364), .B1(new_n463), .B2(new_n467), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n454), .C2(new_n443), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n438), .A2(new_n442), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n289), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n454), .A2(new_n304), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n468), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n468), .ZN(new_n479));
  OAI21_X1  g0279(.A(G200), .B1(new_n443), .B2(new_n454), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n449), .A2(new_n453), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n479), .B(new_n480), .C1(new_n482), .C2(new_n321), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n474), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n283), .A2(new_n209), .A3(G68), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT19), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT81), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT80), .A3(new_n209), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT80), .B1(new_n491), .B2(new_n209), .ZN(new_n494));
  NOR3_X1   g0294(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n247), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n350), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n466), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n349), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n249), .A2(new_n459), .ZN(new_n503));
  AND2_X1   g0303(.A1(G244), .A2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n283), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n373), .A2(new_n375), .A3(G238), .A4(new_n284), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n433), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G250), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n450), .B1(new_n445), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n274), .A3(new_n277), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n304), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n364), .B1(new_n507), .B2(new_n511), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n502), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n486), .A2(new_n487), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n487), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n491), .A2(new_n209), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n495), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n492), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(new_n526), .A3(new_n485), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n500), .B1(new_n527), .B2(new_n247), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n466), .A2(G87), .ZN(new_n529));
  OAI21_X1  g0329(.A(G200), .B1(new_n507), .B2(new_n511), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n373), .A2(new_n375), .A3(new_n504), .ZN(new_n531));
  INV_X1    g0331(.A(new_n503), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n506), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n289), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(G190), .A3(new_n510), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n515), .A2(new_n516), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n516), .B1(new_n515), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n448), .A2(new_n274), .A3(G257), .A4(new_n277), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n453), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n373), .A2(new_n375), .A3(G244), .A4(new_n284), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n284), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n373), .A2(new_n375), .A3(G250), .A4(G1698), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n456), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n541), .B1(new_n547), .B2(new_n289), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n304), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n456), .B(new_n546), .C1(new_n542), .C2(new_n543), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n542), .A2(new_n543), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n289), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n541), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n364), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n253), .A2(G77), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n358), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  XNOR2_X1  g0357(.A(G97), .B(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(new_n209), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT7), .B1(new_n376), .B2(new_n209), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n371), .B(G20), .C1(new_n373), .C2(new_n375), .ZN(new_n563));
  OAI21_X1  g0363(.A(G107), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(KEYINPUT79), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n358), .B1(new_n372), .B2(new_n377), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n354), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n349), .A2(G97), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n466), .B2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n549), .B(new_n555), .C1(new_n569), .C2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n448), .A2(new_n274), .A3(new_n277), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n373), .A2(new_n375), .A3(G257), .A4(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n373), .A2(new_n375), .A3(G250), .A4(new_n284), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n576), .C1(new_n249), .C2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(G264), .A2(new_n574), .B1(new_n578), .B2(new_n289), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n304), .A3(new_n453), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n289), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n448), .A2(new_n274), .A3(G264), .A4(new_n277), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n453), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n364), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n373), .A2(new_n375), .A3(new_n209), .A4(G87), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT22), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n283), .A2(new_n587), .A3(new_n209), .A4(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n209), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n358), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n591), .A2(new_n592), .B1(new_n503), .B2(new_n209), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n354), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n358), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT85), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT25), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n349), .B2(G107), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n466), .A2(G107), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n580), .B(new_n584), .C1(new_n598), .C2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n557), .ZN(new_n609));
  AND2_X1   g0409(.A1(G97), .A2(G107), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n559), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n566), .B2(new_n567), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT79), .B(new_n358), .C1(new_n372), .C2(new_n377), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n247), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n552), .A2(new_n553), .A3(new_n321), .ZN(new_n618));
  AOI21_X1  g0418(.A(G200), .B1(new_n552), .B2(new_n553), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n617), .B(new_n571), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n597), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n596), .B1(new_n589), .B2(new_n593), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n247), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n603), .A2(new_n604), .B1(G107), .B2(new_n466), .ZN(new_n624));
  AOI21_X1  g0424(.A(G200), .B1(new_n579), .B2(new_n453), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n583), .A2(G190), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n573), .A2(new_n608), .A3(new_n620), .A4(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n432), .A2(new_n484), .A3(new_n539), .A4(new_n628), .ZN(G372));
  NAND3_X1  g0429(.A1(new_n474), .A2(new_n478), .A3(new_n608), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n528), .A2(new_n499), .B1(new_n304), .B2(new_n512), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT86), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n509), .A2(new_n633), .A3(new_n274), .A4(new_n277), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n534), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n364), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(KEYINPUT87), .A3(new_n364), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n631), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n635), .A2(G200), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n528), .A3(new_n529), .A4(new_n535), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n640), .A2(new_n627), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n573), .A2(new_n630), .A3(new_n643), .A4(new_n620), .ZN(new_n644));
  INV_X1    g0444(.A(new_n573), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n640), .A4(new_n642), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n537), .A2(new_n538), .A3(new_n573), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n647), .B(new_n640), .C1(new_n648), .C2(new_n646), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n432), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n420), .A2(new_n430), .ZN(new_n651));
  INV_X1    g0451(.A(new_n347), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n367), .A2(KEYINPUT88), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n367), .A2(KEYINPUT88), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n339), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n426), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n300), .A2(new_n301), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n305), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n650), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT89), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G213), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n468), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n484), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n474), .A2(new_n478), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n670), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n669), .B1(new_n598), .B2(new_n607), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n608), .A3(new_n627), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n608), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n669), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT91), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n672), .A2(new_n669), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n669), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n212), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n525), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n228), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n689), .B1(new_n644), .B2(new_n649), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT94), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(KEYINPUT94), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n645), .A2(KEYINPUT26), .A3(new_n640), .A4(new_n642), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n648), .B2(KEYINPUT26), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT95), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n573), .A2(new_n707), .A3(new_n620), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n573), .B2(new_n620), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n630), .B(new_n643), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n710), .A3(new_n640), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n689), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n476), .A2(new_n548), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n579), .A2(new_n477), .A3(new_n512), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT92), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n581), .A2(new_n534), .A3(new_n510), .A4(new_n582), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n481), .A2(G179), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n476), .A4(new_n548), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n635), .A2(new_n304), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n548), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n482), .A3(new_n726), .A4(new_n583), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n554), .A2(new_n304), .A3(new_n583), .A4(new_n635), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT93), .B1(new_n728), .B2(new_n455), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n548), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n669), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n484), .A2(new_n628), .A3(new_n539), .A4(new_n689), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n730), .B1(new_n455), .B2(new_n728), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT31), .B(new_n669), .C1(new_n723), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n713), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT96), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n713), .A2(KEYINPUT96), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n699), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n263), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n208), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n694), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n674), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(new_n304), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n756), .A2(new_n321), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n321), .A2(new_n293), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n209), .A2(G179), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n380), .B1(new_n404), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n755), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G50), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n760), .A2(new_n321), .A3(G200), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G107), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n765), .B(new_n768), .C1(new_n205), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n756), .A2(new_n293), .A3(G190), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n376), .B1(new_n775), .B2(G68), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n760), .A2(new_n769), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT32), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OR3_X1    g0579(.A1(new_n777), .A2(KEYINPUT32), .A3(new_n778), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n321), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n209), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n779), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n775), .A2(new_n786), .B1(new_n757), .B2(G322), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n376), .B1(new_n770), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G294), .B2(new_n783), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT100), .B(G326), .ZN(new_n791));
  INV_X1    g0591(.A(new_n777), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n764), .A2(new_n791), .B1(new_n792), .B2(G329), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n767), .A2(G283), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n761), .B(KEYINPUT101), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n774), .A2(new_n785), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n224), .B1(G20), .B2(new_n364), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n753), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n212), .A2(new_n283), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(KEYINPUT97), .B2(G355), .ZN(new_n804));
  OR2_X1    g0604(.A1(G355), .A2(KEYINPUT97), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(new_n459), .B2(new_n693), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n693), .A2(new_n283), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n227), .A2(new_n444), .A3(G50), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n244), .C2(new_n444), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n750), .B1(new_n754), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n674), .A2(new_n675), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n677), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n750), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT102), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n669), .A2(new_n355), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n369), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n653), .A2(new_n355), .A3(new_n654), .A4(new_n669), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n701), .A2(new_n703), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n689), .C1(new_n644), .C2(new_n649), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n749), .B1(new_n825), .B2(new_n739), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n739), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n801), .A2(new_n751), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n750), .B1(new_n205), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n767), .A2(G87), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n788), .B2(new_n777), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT103), .Z(new_n832));
  INV_X1    g0632(.A(new_n775), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(new_n763), .B2(new_n798), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n283), .B(new_n835), .C1(G294), .C2(new_n757), .ZN(new_n836));
  INV_X1    g0636(.A(new_n773), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G116), .B1(new_n796), .B2(G107), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n784), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT104), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n757), .A2(G143), .B1(new_n764), .B2(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n255), .B2(new_n833), .C1(new_n773), .C2(new_n778), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n796), .A2(G50), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n767), .A2(G68), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n783), .A2(G58), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n376), .B1(new_n792), .B2(G132), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n842), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(KEYINPUT34), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n840), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(KEYINPUT105), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n801), .B1(new_n852), .B2(KEYINPUT105), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n829), .B1(new_n752), .B2(new_n820), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n827), .A2(new_n855), .ZN(G384));
  AND2_X1   g0656(.A1(new_n613), .A2(KEYINPUT35), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n613), .A2(KEYINPUT35), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(new_n459), .A4(new_n226), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n205), .B(new_n228), .C1(new_n308), .C2(G58), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n861), .A2(KEYINPUT106), .B1(G68), .B2(new_n201), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(KEYINPUT106), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n208), .A2(G13), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n432), .A2(new_n704), .A3(new_n712), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n659), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT108), .ZN(new_n868));
  INV_X1    g0668(.A(new_n667), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n426), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n422), .A2(new_n869), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n379), .A2(new_n382), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n384), .B1(KEYINPUT16), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n393), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n874), .B2(new_n429), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n394), .B1(new_n422), .B2(new_n869), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n418), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(KEYINPUT37), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n667), .B1(new_n873), .B2(new_n393), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n431), .A2(KEYINPUT107), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT107), .B1(new_n431), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT38), .B(new_n878), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n346), .A2(new_n669), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n347), .A2(new_n339), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n333), .A2(new_n338), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n346), .B(new_n669), .C1(new_n889), .C2(new_n345), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n367), .A2(new_n669), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n823), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n870), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n431), .A2(new_n394), .A3(new_n869), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n877), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n883), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n347), .A2(new_n669), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n894), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n868), .B(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n891), .A2(new_n821), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT31), .B(new_n669), .C1(new_n723), .C2(new_n731), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n734), .A2(new_n735), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n884), .B2(new_n885), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n914), .B1(new_n900), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n432), .A2(new_n910), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n675), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n919), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n920), .B1(new_n208), .B2(new_n746), .C1(new_n907), .C2(new_n919), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT109), .B1(new_n907), .B2(new_n919), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n865), .B1(new_n921), .B2(new_n922), .ZN(G367));
  INV_X1    g0723(.A(new_n686), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n669), .B1(new_n569), .B2(new_n572), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n708), .B2(new_n709), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n645), .A2(new_n669), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n691), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n691), .A2(new_n929), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n686), .A2(new_n931), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n677), .A2(KEYINPUT112), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n684), .A2(new_n687), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT112), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n688), .C1(new_n676), .C2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n939), .B(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n938), .A2(new_n943), .B1(new_n742), .B2(new_n743), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n694), .B(KEYINPUT41), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n747), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n928), .B(KEYINPUT111), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n682), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n669), .B1(new_n948), .B2(new_n573), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n688), .A2(new_n929), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n528), .A2(new_n529), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n669), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT110), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n640), .A2(new_n642), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n640), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n958), .B2(new_n955), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n950), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT43), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n950), .A2(new_n963), .A3(new_n959), .A4(new_n952), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n947), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n924), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n965), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n946), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n959), .A2(new_n753), .ZN(new_n970));
  INV_X1    g0770(.A(new_n807), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n802), .B1(new_n212), .B2(new_n350), .C1(new_n971), .C2(new_n237), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n749), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n833), .A2(new_n778), .B1(new_n205), .B2(new_n766), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n376), .B(new_n974), .C1(G150), .C2(new_n757), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n783), .A2(G68), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n773), .A2(new_n201), .ZN(new_n977));
  INV_X1    g0777(.A(G143), .ZN(new_n978));
  INV_X1    g0778(.A(G137), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n763), .A2(new_n978), .B1(new_n777), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n761), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(G58), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n283), .B1(new_n775), .B2(G294), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n761), .A2(new_n459), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(KEYINPUT46), .B2(new_n985), .C1(new_n358), .C2(new_n782), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n837), .A2(G283), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n757), .A2(new_n439), .B1(G317), .B2(new_n792), .ZN(new_n989));
  INV_X1    g0789(.A(new_n766), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G311), .A2(new_n764), .B1(new_n990), .B2(G97), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n973), .B1(new_n995), .B2(new_n801), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n970), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n969), .A2(new_n997), .ZN(G387));
  NOR2_X1   g0798(.A1(new_n234), .A2(new_n444), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT114), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n352), .A2(new_n266), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n696), .B(new_n444), .C1(new_n317), .C2(new_n205), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n807), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n999), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(G107), .B2(new_n212), .C1(new_n696), .C2(new_n803), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n750), .B1(new_n1007), .B2(new_n802), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n775), .A2(new_n352), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n783), .A2(new_n498), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n376), .B1(new_n792), .B2(G150), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n981), .A2(G77), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n757), .A2(G50), .B1(new_n764), .B2(G159), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n317), .B2(new_n770), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G97), .C2(new_n767), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n376), .B1(new_n766), .B2(new_n459), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n775), .B1(new_n757), .B2(G317), .ZN(new_n1018));
  INV_X1    g0818(.A(G322), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n763), .C1(new_n773), .C2(new_n436), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n783), .A2(G283), .B1(new_n981), .B2(G294), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT49), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1017), .B(new_n1027), .C1(new_n792), .C2(new_n791), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1016), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n801), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1008), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n684), .B2(new_n753), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n943), .B2(new_n748), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n744), .A2(new_n943), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n694), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n744), .A2(new_n943), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  AND2_X1   g0838(.A1(new_n744), .A2(new_n943), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n695), .B1(new_n1039), .B2(new_n938), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n938), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n1035), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n966), .A2(new_n753), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n802), .B1(new_n457), .B2(new_n212), .C1(new_n971), .C2(new_n241), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n749), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n833), .A2(new_n201), .B1(new_n978), .B2(new_n777), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n376), .B(new_n1047), .C1(new_n308), .C2(new_n981), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n782), .A2(new_n205), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n837), .A2(new_n352), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n830), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n757), .A2(G159), .B1(new_n764), .B2(G150), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n376), .B1(new_n577), .B2(new_n770), .C1(new_n833), .C2(new_n436), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G116), .B2(new_n783), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n757), .A2(G311), .B1(new_n764), .B2(G317), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n761), .A2(new_n834), .B1(new_n777), .B2(new_n1019), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n768), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1052), .A2(new_n1054), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1046), .B1(new_n1064), .B2(new_n801), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n938), .A2(new_n748), .B1(new_n1044), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1043), .A2(new_n1066), .ZN(G390));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n711), .A2(new_n689), .A3(new_n820), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n892), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n892), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n910), .A2(G330), .A3(new_n820), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n891), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n888), .A2(new_n890), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(G330), .A3(new_n738), .A4(new_n820), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1069), .A2(new_n892), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT116), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n892), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n823), .A2(new_n892), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n891), .B1(new_n739), .B2(new_n821), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n908), .A2(G330), .A3(new_n910), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT117), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n891), .C1(new_n739), .C2(new_n821), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1078), .A2(new_n1085), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n432), .A2(G330), .A3(new_n910), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n866), .A2(new_n1094), .A3(new_n659), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT119), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1086), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1072), .A2(new_n1068), .A3(new_n1077), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT118), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT119), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n866), .A2(new_n1094), .A3(new_n659), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n893), .A2(new_n904), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT39), .B1(new_n885), .B2(new_n899), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1081), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n900), .A2(new_n1110), .A3(new_n905), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1111), .A3(new_n1076), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1089), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1105), .B1(new_n895), .B2(new_n902), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1111), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n695), .B1(new_n1104), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT120), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1104), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1089), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1076), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1114), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1118), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n748), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n903), .A2(new_n751), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n828), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n749), .B1(new_n352), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n764), .A2(G128), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n833), .B2(new_n979), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G132), .B2(new_n757), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n981), .A2(G150), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT53), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1135), .A2(KEYINPUT53), .B1(new_n783), .B2(G159), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  NAND2_X1  g0938(.A1(new_n837), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n283), .B1(new_n777), .B2(new_n1141), .C1(new_n201), .C2(new_n766), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT121), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n283), .B(new_n1049), .C1(G283), .C2(new_n764), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G107), .A2(new_n775), .B1(new_n757), .B2(G116), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n577), .C2(new_n777), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n846), .B1(new_n457), .B2(new_n773), .C1(new_n797), .C2(new_n404), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1140), .A2(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1131), .B1(new_n1148), .B2(new_n801), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1129), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1127), .A2(new_n1128), .A3(new_n1150), .ZN(G378));
  AOI22_X1  g0951(.A1(new_n757), .A2(G128), .B1(new_n764), .B2(G125), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n979), .B2(new_n770), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n775), .A2(G132), .B1(new_n981), .B2(new_n1138), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n255), .B2(new_n782), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n792), .A2(G124), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n990), .C2(G159), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n775), .A2(G97), .B1(new_n764), .B2(G116), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n283), .A2(G41), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1163), .A2(new_n1012), .A3(new_n976), .A4(new_n1164), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n380), .A2(new_n766), .B1(new_n770), .B2(new_n350), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n758), .A2(new_n358), .B1(new_n777), .B2(new_n834), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT58), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(KEYINPUT58), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1164), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n266), .C1(G33), .C2(G41), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1162), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n801), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n750), .B1(new_n201), .B2(new_n828), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n296), .A2(new_n869), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT122), .Z(new_n1177));
  XNOR2_X1  g0977(.A(new_n306), .B(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1179));
  XOR2_X1   g0979(.A(new_n1178), .B(new_n1179), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1174), .B(new_n1175), .C1(new_n1181), .C2(new_n752), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n915), .A2(new_n900), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n1183), .C1(new_n912), .C2(KEYINPUT40), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n906), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1184), .B(new_n894), .C1(new_n903), .C2(new_n905), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1180), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1182), .B1(new_n1191), .B2(new_n747), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1102), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1191), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1119), .B1(new_n1104), .B2(new_n1117), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1124), .A2(KEYINPUT120), .A3(new_n1125), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1095), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n694), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1193), .B1(new_n1196), .B2(new_n1201), .ZN(G375));
  INV_X1    g1002(.A(new_n945), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1104), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n891), .A2(new_n751), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n749), .B1(G68), .B2(new_n1130), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n796), .A2(G97), .B1(new_n767), .B2(G77), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n358), .B2(new_n773), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G116), .A2(new_n775), .B1(new_n757), .B2(G283), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n283), .B1(new_n764), .B2(G294), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n792), .A2(G303), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1010), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n764), .A2(G132), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1138), .A2(new_n775), .B1(new_n757), .B2(G137), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n797), .C2(new_n778), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n770), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G150), .A2(new_n1217), .B1(new_n792), .B2(G128), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n376), .B1(new_n990), .B2(G58), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n266), .C2(new_n782), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1209), .A2(new_n1213), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1207), .B1(new_n1221), .B2(new_n801), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1100), .A2(new_n748), .B1(new_n1206), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1205), .A2(new_n1223), .ZN(G381));
  INV_X1    g1024(.A(new_n1200), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n695), .B1(new_n1225), .B2(new_n1194), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1199), .B2(new_n1191), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1192), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G390), .ZN(new_n1230));
  INV_X1    g1030(.A(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1232), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1127), .A2(new_n1128), .A3(new_n1150), .ZN(new_n1234));
  INV_X1    g1034(.A(G381), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1229), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT123), .Z(G407));
  NAND3_X1  g1037(.A1(new_n1229), .A2(new_n668), .A3(new_n1234), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  OAI211_X1 g1039(.A(G378), .B(new_n1193), .C1(new_n1196), .C2(new_n1201), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1199), .A2(new_n945), .A3(new_n1191), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1241), .B2(new_n1192), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1204), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n694), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1104), .A2(new_n1204), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(KEYINPUT60), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(G384), .A3(new_n1223), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1223), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1231), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G213), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(G343), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1243), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(KEYINPUT126), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(G2897), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1253), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1250), .A2(new_n1252), .A3(new_n1263), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1194), .A2(new_n1203), .A3(new_n1195), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G378), .B1(new_n1268), .B2(new_n1193), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1229), .B2(G378), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1270), .B2(new_n1256), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1256), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1254), .A3(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1261), .A2(new_n1262), .A3(new_n1271), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1230), .ZN(new_n1276));
  XOR2_X1   g1076(.A(G393), .B(G396), .Z(new_n1277));
  AOI22_X1  g1077(.A1(new_n946), .A2(new_n968), .B1(new_n970), .B2(new_n996), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(G390), .ZN(new_n1279));
  AND4_X1   g1079(.A1(KEYINPUT124), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1278), .B2(G390), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1282), .A2(new_n1277), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT127), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1275), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1254), .A4(new_n1257), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT125), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1272), .A2(new_n1289), .A3(KEYINPUT63), .A4(new_n1254), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1262), .B(new_n1292), .C1(new_n1272), .C2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1254), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1286), .A2(new_n1297), .ZN(G405));
  NAND2_X1  g1098(.A1(G375), .A2(new_n1234), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1240), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1254), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1253), .A3(new_n1240), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1284), .ZN(G402));
endmodule


