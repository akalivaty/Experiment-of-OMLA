

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753;

  AND2_X1 U366 ( .A1(n392), .A2(n390), .ZN(n389) );
  NOR2_X1 U367 ( .A1(n520), .A2(n519), .ZN(n642) );
  XNOR2_X1 U368 ( .A(n526), .B(KEYINPUT33), .ZN(n413) );
  BUF_X1 U369 ( .A(n698), .Z(n347) );
  XNOR2_X1 U370 ( .A(n524), .B(KEYINPUT78), .ZN(n535) );
  XNOR2_X1 U371 ( .A(n579), .B(KEYINPUT1), .ZN(n698) );
  OR2_X1 U372 ( .A1(n673), .A2(G902), .ZN(n364) );
  XNOR2_X1 U373 ( .A(n501), .B(n500), .ZN(n673) );
  XNOR2_X1 U374 ( .A(n424), .B(n494), .ZN(n394) );
  AND2_X2 U375 ( .A1(n412), .A2(n357), .ZN(n363) );
  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U377 ( .A(G137), .B(G128), .ZN(n378) );
  NAND2_X1 U378 ( .A1(n581), .A2(n447), .ZN(n350) );
  NAND2_X1 U379 ( .A1(n552), .A2(n551), .ZN(n348) );
  XNOR2_X2 U380 ( .A(n485), .B(n484), .ZN(n552) );
  XNOR2_X2 U381 ( .A(n452), .B(n451), .ZN(n487) );
  XNOR2_X2 U382 ( .A(n498), .B(n497), .ZN(n704) );
  INV_X1 U383 ( .A(n647), .ZN(n503) );
  INV_X1 U384 ( .A(KEYINPUT74), .ZN(n409) );
  INV_X2 U385 ( .A(G953), .ZN(n650) );
  NOR2_X1 U386 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U387 ( .A1(n361), .A2(n359), .ZN(n485) );
  OR2_X1 U388 ( .A1(n543), .A2(n538), .ZN(n714) );
  XNOR2_X1 U389 ( .A(n737), .B(n409), .ZN(n425) );
  INV_X1 U390 ( .A(n448), .ZN(n349) );
  XNOR2_X1 U391 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n428) );
  XNOR2_X1 U392 ( .A(G125), .B(G146), .ZN(n465) );
  INV_X1 U393 ( .A(n361), .ZN(n527) );
  XNOR2_X2 U394 ( .A(n350), .B(n349), .ZN(n361) );
  XNOR2_X2 U395 ( .A(n570), .B(n440), .ZN(n581) );
  NOR2_X2 U396 ( .A1(n660), .A2(n642), .ZN(n521) );
  XNOR2_X1 U397 ( .A(n407), .B(n355), .ZN(n404) );
  NOR2_X1 U398 ( .A1(n645), .A2(n391), .ZN(n390) );
  INV_X1 U399 ( .A(KEYINPUT84), .ZN(n419) );
  OR2_X1 U400 ( .A1(n704), .A2(n611), .ZN(n589) );
  AND2_X1 U401 ( .A1(n406), .A2(n600), .ZN(n401) );
  AND2_X1 U402 ( .A1(n406), .A2(n381), .ZN(n399) );
  XNOR2_X1 U403 ( .A(n486), .B(G137), .ZN(n414) );
  INV_X1 U404 ( .A(n634), .ZN(n362) );
  INV_X1 U405 ( .A(n663), .ZN(n496) );
  XNOR2_X1 U406 ( .A(n482), .B(n360), .ZN(n359) );
  INV_X1 U407 ( .A(KEYINPUT104), .ZN(n360) );
  BUF_X1 U408 ( .A(n522), .Z(n566) );
  NAND2_X1 U409 ( .A1(n366), .A2(n411), .ZN(n365) );
  XNOR2_X1 U410 ( .A(n537), .B(n372), .ZN(n544) );
  INV_X1 U411 ( .A(KEYINPUT31), .ZN(n372) );
  XNOR2_X1 U412 ( .A(n659), .B(n575), .ZN(n406) );
  INV_X1 U413 ( .A(G237), .ZN(n434) );
  NOR2_X1 U414 ( .A1(n662), .A2(KEYINPUT70), .ZN(n534) );
  INV_X1 U415 ( .A(KEYINPUT44), .ZN(n386) );
  XNOR2_X1 U416 ( .A(n464), .B(n465), .ZN(n647) );
  XNOR2_X1 U417 ( .A(n398), .B(KEYINPUT98), .ZN(n397) );
  XNOR2_X1 U418 ( .A(G113), .B(G122), .ZN(n467) );
  XNOR2_X1 U419 ( .A(n394), .B(n425), .ZN(n433) );
  NAND2_X1 U420 ( .A1(G237), .A2(G234), .ZN(n441) );
  XNOR2_X1 U421 ( .A(n704), .B(KEYINPUT6), .ZN(n567) );
  XNOR2_X1 U422 ( .A(n501), .B(n353), .ZN(n663) );
  NAND2_X1 U423 ( .A1(n620), .A2(n619), .ZN(n646) );
  INV_X1 U424 ( .A(KEYINPUT24), .ZN(n380) );
  XNOR2_X1 U425 ( .A(G119), .B(KEYINPUT23), .ZN(n376) );
  XNOR2_X1 U426 ( .A(G110), .B(KEYINPUT92), .ZN(n375) );
  INV_X1 U427 ( .A(G134), .ZN(n451) );
  XNOR2_X1 U428 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n454) );
  XOR2_X1 U429 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n455) );
  INV_X1 U430 ( .A(KEYINPUT41), .ZN(n607) );
  XNOR2_X1 U431 ( .A(n477), .B(n476), .ZN(n538) );
  AND2_X1 U432 ( .A1(n593), .A2(n592), .ZN(n602) );
  NAND2_X1 U433 ( .A1(n370), .A2(n368), .ZN(n384) );
  NAND2_X1 U434 ( .A1(n369), .A2(n411), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n425), .B(n352), .ZN(n500) );
  INV_X1 U436 ( .A(G104), .ZN(n640) );
  XNOR2_X1 U437 ( .A(n556), .B(KEYINPUT106), .ZN(n645) );
  AND2_X1 U438 ( .A1(n544), .A2(n371), .ZN(n695) );
  INV_X1 U439 ( .A(n694), .ZN(n371) );
  AND2_X1 U440 ( .A1(n544), .A2(n373), .ZN(n644) );
  AND2_X1 U441 ( .A1(n609), .A2(n354), .ZN(n351) );
  XOR2_X1 U442 ( .A(n499), .B(G140), .Z(n352) );
  XOR2_X1 U443 ( .A(n495), .B(n494), .Z(n353) );
  AND2_X2 U444 ( .A1(n384), .A2(n626), .ZN(n678) );
  AND2_X1 U445 ( .A1(n582), .A2(n373), .ZN(n354) );
  XOR2_X1 U446 ( .A(KEYINPUT86), .B(KEYINPUT46), .Z(n355) );
  XNOR2_X1 U447 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n356) );
  INV_X1 U448 ( .A(KEYINPUT65), .ZN(n411) );
  AND2_X1 U449 ( .A1(n624), .A2(KEYINPUT65), .ZN(n357) );
  NAND2_X1 U450 ( .A1(KEYINPUT84), .A2(n621), .ZN(n358) );
  INV_X1 U451 ( .A(KEYINPUT48), .ZN(n405) );
  NAND2_X1 U452 ( .A1(n525), .A2(n567), .ZN(n526) );
  NAND2_X1 U453 ( .A1(n362), .A2(n507), .ZN(n477) );
  NAND2_X1 U454 ( .A1(n396), .A2(n363), .ZN(n367) );
  NAND2_X1 U455 ( .A1(n496), .A2(n507), .ZN(n498) );
  XNOR2_X2 U456 ( .A(n649), .B(n489), .ZN(n501) );
  XNOR2_X2 U457 ( .A(n364), .B(G469), .ZN(n579) );
  AND2_X2 U458 ( .A1(n367), .A2(n365), .ZN(n370) );
  NAND2_X1 U459 ( .A1(n412), .A2(n624), .ZN(n366) );
  INV_X1 U460 ( .A(n396), .ZN(n369) );
  NAND2_X1 U461 ( .A1(n609), .A2(n582), .ZN(n374) );
  INV_X1 U462 ( .A(n643), .ZN(n373) );
  NOR2_X1 U463 ( .A1(n374), .A2(n694), .ZN(n692) );
  NOR2_X1 U464 ( .A1(n584), .A2(n374), .ZN(n585) );
  XNOR2_X1 U465 ( .A(n376), .B(n375), .ZN(n379) );
  XNOR2_X1 U466 ( .A(n379), .B(n377), .ZN(n502) );
  XNOR2_X1 U467 ( .A(n378), .B(n380), .ZN(n377) );
  AND2_X1 U468 ( .A1(n600), .A2(KEYINPUT48), .ZN(n381) );
  NAND2_X1 U469 ( .A1(n574), .A2(n347), .ZN(n659) );
  INV_X1 U470 ( .A(n535), .ZN(n525) );
  NAND2_X2 U471 ( .A1(n382), .A2(n383), .ZN(n570) );
  INV_X1 U472 ( .A(n594), .ZN(n382) );
  XNOR2_X1 U473 ( .A(n437), .B(n436), .ZN(n594) );
  INV_X1 U474 ( .A(n611), .ZN(n383) );
  NAND2_X1 U475 ( .A1(n389), .A2(n385), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n387), .B(n386), .ZN(n385) );
  NAND2_X1 U477 ( .A1(n388), .A2(n662), .ZN(n387) );
  XNOR2_X2 U478 ( .A(n533), .B(n532), .ZN(n662) );
  NOR2_X1 U479 ( .A1(n558), .A2(n557), .ZN(n388) );
  NAND2_X1 U480 ( .A1(n550), .A2(n549), .ZN(n391) );
  NAND2_X1 U481 ( .A1(n393), .A2(n534), .ZN(n392) );
  INV_X1 U482 ( .A(n558), .ZN(n393) );
  XNOR2_X1 U483 ( .A(n738), .B(n394), .ZN(n740) );
  AND2_X1 U484 ( .A1(n417), .A2(n395), .ZN(n625) );
  INV_X1 U485 ( .A(n646), .ZN(n395) );
  AND2_X1 U486 ( .A1(n417), .A2(n650), .ZN(n741) );
  XNOR2_X2 U487 ( .A(n410), .B(n356), .ZN(n417) );
  NAND2_X1 U488 ( .A1(n415), .A2(n419), .ZN(n396) );
  XNOR2_X1 U489 ( .A(n397), .B(n486), .ZN(n466) );
  NAND2_X1 U490 ( .A1(n490), .A2(G214), .ZN(n398) );
  NAND2_X1 U491 ( .A1(n399), .A2(n404), .ZN(n402) );
  NAND2_X1 U492 ( .A1(n400), .A2(n405), .ZN(n403) );
  NAND2_X1 U493 ( .A1(n401), .A2(n404), .ZN(n400) );
  NAND2_X1 U494 ( .A1(n403), .A2(n402), .ZN(n620) );
  NAND2_X1 U495 ( .A1(n751), .A2(n752), .ZN(n407) );
  INV_X1 U496 ( .A(n538), .ZN(n542) );
  XNOR2_X2 U497 ( .A(n408), .B(KEYINPUT102), .ZN(n643) );
  NAND2_X1 U498 ( .A1(n539), .A2(n538), .ZN(n408) );
  NAND2_X1 U499 ( .A1(n418), .A2(n417), .ZN(n412) );
  NAND2_X1 U500 ( .A1(n413), .A2(n547), .ZN(n529) );
  NAND2_X1 U501 ( .A1(n413), .A2(n722), .ZN(n723) );
  AND2_X1 U502 ( .A1(n413), .A2(n729), .ZN(n730) );
  XNOR2_X2 U503 ( .A(n487), .B(n414), .ZN(n649) );
  NAND2_X1 U504 ( .A1(n417), .A2(n416), .ZN(n415) );
  NOR2_X1 U505 ( .A1(n646), .A2(n623), .ZN(n416) );
  NOR2_X1 U506 ( .A1(n646), .A2(n358), .ZN(n418) );
  BUF_X1 U507 ( .A(n660), .Z(n661) );
  XNOR2_X1 U508 ( .A(n516), .B(n515), .ZN(n660) );
  XNOR2_X1 U509 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n420) );
  INV_X1 U510 ( .A(KEYINPUT70), .ZN(n557) );
  INV_X1 U511 ( .A(KEYINPUT87), .ZN(n575) );
  INV_X1 U512 ( .A(KEYINPUT124), .ZN(n631) );
  XNOR2_X1 U513 ( .A(n605), .B(n420), .ZN(n751) );
  XNOR2_X2 U514 ( .A(G110), .B(G107), .ZN(n421) );
  XNOR2_X2 U515 ( .A(n421), .B(G104), .ZN(n737) );
  XNOR2_X2 U516 ( .A(KEYINPUT3), .B(G119), .ZN(n422) );
  XNOR2_X2 U517 ( .A(n422), .B(G113), .ZN(n494) );
  XNOR2_X2 U518 ( .A(G122), .B(G116), .ZN(n456) );
  XNOR2_X1 U519 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n423) );
  XNOR2_X1 U520 ( .A(n456), .B(n423), .ZN(n424) );
  XNOR2_X1 U521 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U522 ( .A(n426), .B(G101), .ZN(n488) );
  NAND2_X1 U523 ( .A1(n650), .A2(G224), .ZN(n427) );
  XNOR2_X1 U524 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n488), .B(n429), .ZN(n431) );
  XNOR2_X2 U526 ( .A(G143), .B(G128), .ZN(n452) );
  XNOR2_X1 U527 ( .A(n452), .B(n465), .ZN(n430) );
  XNOR2_X1 U528 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U529 ( .A(n433), .B(n432), .ZN(n679) );
  XNOR2_X1 U530 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  INV_X1 U531 ( .A(n623), .ZN(n621) );
  NOR2_X1 U532 ( .A1(n679), .A2(n621), .ZN(n437) );
  INV_X1 U533 ( .A(G902), .ZN(n507) );
  NAND2_X1 U534 ( .A1(n507), .A2(n434), .ZN(n438) );
  NAND2_X1 U535 ( .A1(n438), .A2(G210), .ZN(n435) );
  XOR2_X1 U536 ( .A(n435), .B(KEYINPUT90), .Z(n436) );
  AND2_X1 U537 ( .A1(n438), .A2(G214), .ZN(n611) );
  INV_X1 U538 ( .A(KEYINPUT79), .ZN(n439) );
  XNOR2_X1 U539 ( .A(n439), .B(KEYINPUT19), .ZN(n440) );
  XOR2_X1 U540 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n442) );
  XNOR2_X1 U541 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U542 ( .A1(G952), .A2(n443), .ZN(n727) );
  OR2_X1 U543 ( .A1(n727), .A2(G953), .ZN(n562) );
  AND2_X1 U544 ( .A1(G902), .A2(n443), .ZN(n560) );
  INV_X1 U545 ( .A(G898), .ZN(n444) );
  NAND2_X1 U546 ( .A1(n444), .A2(G953), .ZN(n445) );
  XNOR2_X1 U547 ( .A(n445), .B(KEYINPUT91), .ZN(n739) );
  NAND2_X1 U548 ( .A1(n560), .A2(n739), .ZN(n446) );
  NAND2_X1 U549 ( .A1(n562), .A2(n446), .ZN(n447) );
  XNOR2_X1 U550 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n448) );
  XOR2_X1 U551 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n450) );
  NAND2_X1 U552 ( .A1(n650), .A2(G234), .ZN(n449) );
  XNOR2_X1 U553 ( .A(n450), .B(n449), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n504), .A2(G217), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n487), .B(n453), .ZN(n460) );
  XNOR2_X1 U556 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U557 ( .A(n456), .B(G107), .ZN(n457) );
  XNOR2_X1 U558 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n460), .B(n459), .ZN(n670) );
  NAND2_X1 U560 ( .A1(n670), .A2(n507), .ZN(n462) );
  INV_X1 U561 ( .A(G478), .ZN(n461) );
  XNOR2_X1 U562 ( .A(n462), .B(n461), .ZN(n539) );
  INV_X1 U563 ( .A(n539), .ZN(n543) );
  XNOR2_X2 U564 ( .A(KEYINPUT73), .B(G131), .ZN(n486) );
  INV_X1 U565 ( .A(KEYINPUT10), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n463), .B(G140), .ZN(n464) );
  XNOR2_X1 U567 ( .A(n466), .B(n503), .ZN(n474) );
  XNOR2_X1 U568 ( .A(n640), .B(G143), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n468), .B(n467), .ZN(n472) );
  XNOR2_X1 U570 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n470) );
  XNOR2_X1 U571 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U572 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U574 ( .A(n474), .B(n473), .ZN(n634) );
  XNOR2_X1 U575 ( .A(KEYINPUT13), .B(G475), .ZN(n475) );
  XNOR2_X1 U576 ( .A(n475), .B(KEYINPUT99), .ZN(n476) );
  INV_X1 U577 ( .A(n714), .ZN(n481) );
  XOR2_X1 U578 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n480) );
  NAND2_X1 U579 ( .A1(n623), .A2(G234), .ZN(n478) );
  XNOR2_X1 U580 ( .A(n478), .B(KEYINPUT20), .ZN(n508) );
  NAND2_X1 U581 ( .A1(n508), .A2(G221), .ZN(n479) );
  XOR2_X1 U582 ( .A(n480), .B(n479), .Z(n701) );
  NAND2_X1 U583 ( .A1(n481), .A2(n701), .ZN(n482) );
  INV_X1 U584 ( .A(KEYINPUT66), .ZN(n483) );
  XNOR2_X1 U585 ( .A(n483), .B(KEYINPUT22), .ZN(n484) );
  XNOR2_X1 U586 ( .A(n488), .B(G146), .ZN(n489) );
  NAND2_X1 U587 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n491), .B(KEYINPUT5), .ZN(n493) );
  XNOR2_X1 U589 ( .A(G116), .B(KEYINPUT94), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n493), .B(n492), .ZN(n495) );
  INV_X1 U591 ( .A(G472), .ZN(n497) );
  INV_X1 U592 ( .A(n567), .ZN(n551) );
  NAND2_X1 U593 ( .A1(n650), .A2(G227), .ZN(n499) );
  INV_X1 U594 ( .A(n347), .ZN(n553) );
  XNOR2_X1 U595 ( .A(n503), .B(n502), .ZN(n506) );
  NAND2_X1 U596 ( .A1(n504), .A2(G221), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n506), .B(n505), .ZN(n627) );
  NAND2_X1 U598 ( .A1(n627), .A2(n507), .ZN(n512) );
  NAND2_X1 U599 ( .A1(G217), .A2(n508), .ZN(n510) );
  XNOR2_X1 U600 ( .A(KEYINPUT80), .B(KEYINPUT25), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n522) );
  XNOR2_X1 U603 ( .A(n566), .B(KEYINPUT105), .ZN(n702) );
  NOR2_X1 U604 ( .A1(n553), .A2(n702), .ZN(n513) );
  AND2_X1 U605 ( .A1(n551), .A2(n513), .ZN(n514) );
  NAND2_X1 U606 ( .A1(n552), .A2(n514), .ZN(n516) );
  INV_X1 U607 ( .A(KEYINPUT32), .ZN(n515) );
  INV_X1 U608 ( .A(n552), .ZN(n520) );
  INV_X1 U609 ( .A(n704), .ZN(n545) );
  INV_X1 U610 ( .A(n566), .ZN(n517) );
  NOR2_X1 U611 ( .A1(n545), .A2(n517), .ZN(n518) );
  NAND2_X1 U612 ( .A1(n553), .A2(n518), .ZN(n519) );
  XNOR2_X1 U613 ( .A(n521), .B(KEYINPUT89), .ZN(n558) );
  INV_X1 U614 ( .A(n701), .ZN(n564) );
  OR2_X1 U615 ( .A1(n522), .A2(n564), .ZN(n523) );
  XNOR2_X2 U616 ( .A(n523), .B(KEYINPUT71), .ZN(n697) );
  NAND2_X1 U617 ( .A1(n698), .A2(n697), .ZN(n524) );
  INV_X1 U618 ( .A(n527), .ZN(n547) );
  INV_X1 U619 ( .A(KEYINPUT34), .ZN(n528) );
  XNOR2_X1 U620 ( .A(n529), .B(n528), .ZN(n531) );
  OR2_X1 U621 ( .A1(n539), .A2(n542), .ZN(n595) );
  XOR2_X1 U622 ( .A(n595), .B(KEYINPUT82), .Z(n530) );
  NAND2_X1 U623 ( .A1(n531), .A2(n530), .ZN(n533) );
  XNOR2_X1 U624 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n532) );
  NOR2_X1 U625 ( .A1(n535), .A2(n704), .ZN(n536) );
  XNOR2_X1 U626 ( .A(n536), .B(KEYINPUT95), .ZN(n709) );
  NOR2_X1 U627 ( .A1(n709), .A2(n527), .ZN(n537) );
  OR2_X1 U628 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U629 ( .A(KEYINPUT103), .ZN(n540) );
  XNOR2_X1 U630 ( .A(n541), .B(n540), .ZN(n694) );
  NAND2_X1 U631 ( .A1(n694), .A2(n643), .ZN(n718) );
  NAND2_X1 U632 ( .A1(n544), .A2(n718), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n697), .A2(n579), .ZN(n587) );
  NOR2_X1 U634 ( .A1(n587), .A2(n545), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U636 ( .A1(n548), .A2(n694), .ZN(n689) );
  NOR2_X1 U637 ( .A1(n548), .A2(n643), .ZN(n641) );
  NOR2_X1 U638 ( .A1(n689), .A2(n641), .ZN(n549) );
  XNOR2_X1 U639 ( .A(n348), .B(KEYINPUT88), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n553), .A2(n702), .ZN(n554) );
  NOR2_X1 U641 ( .A1(n650), .A2(G900), .ZN(n559) );
  NAND2_X1 U642 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n562), .A2(n561), .ZN(n590) );
  INV_X1 U644 ( .A(n590), .ZN(n563) );
  NOR2_X1 U645 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n566), .A2(n565), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n643), .A2(n576), .ZN(n568) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U649 ( .A(n569), .B(KEYINPUT107), .ZN(n613) );
  XNOR2_X1 U650 ( .A(n613), .B(KEYINPUT113), .ZN(n571) );
  NOR2_X1 U651 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U652 ( .A(KEYINPUT114), .B(KEYINPUT36), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n573), .B(n572), .ZN(n574) );
  OR2_X1 U654 ( .A1(n704), .A2(n576), .ZN(n578) );
  INV_X1 U655 ( .A(KEYINPUT28), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n578), .B(n577), .ZN(n580) );
  AND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n609) );
  BUF_X1 U658 ( .A(n581), .Z(n582) );
  OR2_X1 U659 ( .A1(n351), .A2(KEYINPUT47), .ZN(n583) );
  NOR2_X1 U660 ( .A1(n583), .A2(n692), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n718), .A2(KEYINPUT47), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n599) );
  XNOR2_X1 U663 ( .A(KEYINPUT109), .B(n587), .ZN(n593) );
  INV_X1 U664 ( .A(KEYINPUT30), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n589), .B(n588), .ZN(n591) );
  AND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  BUF_X1 U667 ( .A(n594), .Z(n601) );
  NOR2_X1 U668 ( .A1(n595), .A2(n601), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n602), .A2(n596), .ZN(n597) );
  XNOR2_X1 U670 ( .A(n597), .B(KEYINPUT110), .ZN(n750) );
  XNOR2_X1 U671 ( .A(n750), .B(KEYINPUT83), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT38), .ZN(n713) );
  NAND2_X1 U674 ( .A1(n602), .A2(n713), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n617) );
  NOR2_X1 U677 ( .A1(n617), .A2(n643), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n713), .A2(n383), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT112), .ZN(n717) );
  NOR2_X1 U680 ( .A1(n717), .A2(n714), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(n607), .ZN(n729) );
  NAND2_X1 U682 ( .A1(n729), .A2(n609), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT42), .ZN(n752) );
  NOR2_X1 U684 ( .A1(n347), .A2(n611), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT43), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n615), .A2(n601), .ZN(n616) );
  XOR2_X1 U688 ( .A(KEYINPUT108), .B(n616), .Z(n749) );
  OR2_X1 U689 ( .A1(n617), .A2(n694), .ZN(n696) );
  INV_X1 U690 ( .A(n696), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n749), .A2(n618), .ZN(n619) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n622) );
  OR2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n678), .A2(G217), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n630) );
  INV_X1 U697 ( .A(G952), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n629), .A2(G953), .ZN(n683) );
  NAND2_X1 U699 ( .A1(n630), .A2(n683), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(G66) );
  NAND2_X1 U701 ( .A1(n678), .A2(G475), .ZN(n636) );
  XOR2_X1 U702 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n637), .A2(n683), .ZN(n639) );
  INV_X1 U706 ( .A(KEYINPUT60), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(G60) );
  XOR2_X1 U708 ( .A(G146), .B(n351), .Z(G48) );
  XNOR2_X1 U709 ( .A(n641), .B(n640), .ZN(G6) );
  XOR2_X1 U710 ( .A(G110), .B(n642), .Z(G12) );
  XOR2_X1 U711 ( .A(G113), .B(n644), .Z(G15) );
  XOR2_X1 U712 ( .A(G101), .B(n645), .Z(G3) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT4), .ZN(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n652) );
  XNOR2_X1 U715 ( .A(n646), .B(n652), .ZN(n651) );
  NAND2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n656) );
  XNOR2_X1 U717 ( .A(n652), .B(G227), .ZN(n653) );
  NAND2_X1 U718 ( .A1(n653), .A2(G900), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n654), .A2(G953), .ZN(n655) );
  NAND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(G72) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n657) );
  XOR2_X1 U722 ( .A(n657), .B(G125), .Z(n658) );
  XNOR2_X1 U723 ( .A(n659), .B(n658), .ZN(G27) );
  XOR2_X1 U724 ( .A(n661), .B(G119), .Z(G21) );
  XNOR2_X1 U725 ( .A(n662), .B(G122), .ZN(G24) );
  NAND2_X1 U726 ( .A1(n678), .A2(G472), .ZN(n665) );
  XOR2_X1 U727 ( .A(KEYINPUT62), .B(n663), .Z(n664) );
  XNOR2_X1 U728 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n666), .A2(n683), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n667) );
  XNOR2_X1 U731 ( .A(n668), .B(n667), .ZN(G57) );
  NAND2_X1 U732 ( .A1(n678), .A2(G478), .ZN(n669) );
  XOR2_X1 U733 ( .A(n670), .B(n669), .Z(n671) );
  INV_X1 U734 ( .A(n683), .ZN(n676) );
  NOR2_X1 U735 ( .A1(n671), .A2(n676), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n678), .A2(G469), .ZN(n675) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n672) );
  XNOR2_X1 U738 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(G54) );
  NAND2_X1 U741 ( .A1(n678), .A2(G210), .ZN(n682) );
  XNOR2_X1 U742 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n680) );
  XNOR2_X1 U743 ( .A(n679), .B(n680), .ZN(n681) );
  XNOR2_X1 U744 ( .A(n682), .B(n681), .ZN(n684) );
  NAND2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n687) );
  XOR2_X1 U746 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT85), .ZN(n686) );
  XNOR2_X1 U748 ( .A(n687), .B(n686), .ZN(G51) );
  XNOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n688) );
  XNOR2_X1 U750 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U751 ( .A(G107), .B(n690), .ZN(G9) );
  XNOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n691) );
  XNOR2_X1 U753 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(G128), .B(n693), .ZN(G30) );
  XOR2_X1 U755 ( .A(G116), .B(n695), .Z(G18) );
  XNOR2_X1 U756 ( .A(G134), .B(n696), .ZN(G36) );
  XNOR2_X1 U757 ( .A(n625), .B(KEYINPUT2), .ZN(n734) );
  XNOR2_X1 U758 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n726) );
  NOR2_X1 U759 ( .A1(n347), .A2(n697), .ZN(n700) );
  XOR2_X1 U760 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n699) );
  XNOR2_X1 U761 ( .A(n700), .B(n699), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U763 ( .A(KEYINPUT49), .B(n703), .ZN(n705) );
  AND2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n710), .B(KEYINPUT119), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT51), .ZN(n712) );
  NAND2_X1 U769 ( .A1(n712), .A2(n729), .ZN(n724) );
  NOR2_X1 U770 ( .A1(n713), .A2(n383), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U772 ( .A(KEYINPUT120), .B(n716), .Z(n721) );
  INV_X1 U773 ( .A(n717), .ZN(n719) );
  NAND2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n732), .B(KEYINPUT122), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U782 ( .A1(n735), .A2(G953), .ZN(n736) );
  XNOR2_X1 U783 ( .A(n736), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U784 ( .A(n737), .B(G101), .ZN(n738) );
  OR2_X1 U785 ( .A1(n740), .A2(n739), .ZN(n747) );
  XNOR2_X1 U786 ( .A(n741), .B(KEYINPUT125), .ZN(n745) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(G898), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U791 ( .A(n747), .B(n746), .ZN(n748) );
  XOR2_X1 U792 ( .A(KEYINPUT126), .B(n748), .Z(G69) );
  XOR2_X1 U793 ( .A(G140), .B(n749), .Z(G42) );
  XNOR2_X1 U794 ( .A(G143), .B(n750), .ZN(G45) );
  XNOR2_X1 U795 ( .A(G131), .B(n751), .ZN(G33) );
  XOR2_X1 U796 ( .A(G137), .B(n752), .Z(n753) );
  XNOR2_X1 U797 ( .A(KEYINPUT127), .B(n753), .ZN(G39) );
endmodule

