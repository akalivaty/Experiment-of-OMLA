

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(G160), .A2(G40), .ZN(n705) );
  NOR2_X1 U553 ( .A1(G2105), .A2(n522), .ZN(n597) );
  AND2_X2 U554 ( .A1(n604), .A2(n603), .ZN(n776) );
  INV_X2 U555 ( .A(n657), .ZN(n674) );
  AND2_X4 U556 ( .A1(n704), .A2(n605), .ZN(n657) );
  NOR2_X2 U557 ( .A1(n530), .A2(n529), .ZN(G160) );
  BUF_X2 U558 ( .A(n597), .Z(n909) );
  AND2_X1 U559 ( .A1(n522), .A2(G2105), .ZN(n598) );
  INV_X1 U560 ( .A(G2104), .ZN(n522) );
  NOR2_X1 U561 ( .A1(G543), .A2(n536), .ZN(n531) );
  XNOR2_X1 U562 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X2 U563 ( .A1(G651), .A2(n572), .ZN(n617) );
  XOR2_X2 U564 ( .A(KEYINPUT1), .B(n531), .Z(n634) );
  NOR2_X2 U565 ( .A1(n572), .A2(n536), .ZN(n616) );
  XOR2_X1 U566 ( .A(n615), .B(KEYINPUT31), .Z(n517) );
  OR2_X1 U567 ( .A1(G301), .A2(n669), .ZN(n518) );
  NOR2_X1 U568 ( .A1(n682), .A2(n606), .ZN(n519) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT32), .Z(n520) );
  INV_X1 U570 ( .A(G8), .ZN(n606) );
  NOR2_X1 U571 ( .A1(G1966), .A2(n741), .ZN(n685) );
  XNOR2_X1 U572 ( .A(n681), .B(n520), .ZN(n689) );
  NAND2_X1 U573 ( .A1(G8), .A2(n674), .ZN(n741) );
  INV_X1 U574 ( .A(KEYINPUT103), .ZN(n702) );
  BUF_X2 U575 ( .A(n598), .Z(n902) );
  NOR2_X2 U576 ( .A1(n776), .A2(G1384), .ZN(n704) );
  XOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .Z(n572) );
  INV_X1 U578 ( .A(KEYINPUT71), .ZN(n556) );
  INV_X1 U579 ( .A(KEYINPUT5), .ZN(n539) );
  XNOR2_X1 U580 ( .A(n539), .B(KEYINPUT78), .ZN(n540) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n805) );
  AND2_X2 U582 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  XNOR2_X1 U583 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U584 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NOR2_X2 U585 ( .A1(n638), .A2(n637), .ZN(n937) );
  XOR2_X1 U586 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  NAND2_X1 U587 ( .A1(G101), .A2(n597), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n521), .Z(n525) );
  NAND2_X1 U589 ( .A1(G125), .A2(n598), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n530) );
  NAND2_X1 U591 ( .A1(G113), .A2(n901), .ZN(n528) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT17), .B(n526), .Z(n706) );
  NAND2_X1 U594 ( .A1(G137), .A2(n706), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U596 ( .A1(G51), .A2(n617), .ZN(n533) );
  INV_X1 U597 ( .A(G651), .ZN(n536) );
  NAND2_X1 U598 ( .A1(G63), .A2(n634), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT6), .B(n534), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n805), .A2(G89), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT4), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G76), .A2(n616), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n617), .A2(G52), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(n545), .Z(n547) );
  NAND2_X1 U608 ( .A1(n634), .A2(G64), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(KEYINPUT68), .B(n548), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n805), .A2(G90), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(n549), .Z(n551) );
  NAND2_X1 U613 ( .A1(n616), .A2(G77), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U616 ( .A1(n554), .A2(n553), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(n617), .A2(G53), .ZN(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT72), .B(n555), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n634), .A2(G65), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(n560), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n616), .A2(G78), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G91), .A2(n805), .ZN(n561) );
  AND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(G299) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G75), .A2(n616), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G88), .A2(n805), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G50), .A2(n617), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G62), .A2(n634), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n570), .A2(n569), .ZN(G166) );
  NAND2_X1 U635 ( .A1(G49), .A2(n617), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT82), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G87), .A2(n572), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n634), .A2(n575), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(G288) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  NAND2_X1 U643 ( .A1(n617), .A2(G48), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT86), .B(n578), .ZN(n588) );
  XOR2_X1 U645 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n580) );
  NAND2_X1 U646 ( .A1(G73), .A2(n616), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G86), .A2(n805), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G61), .A2(n634), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT83), .B(n583), .Z(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U653 ( .A(KEYINPUT85), .B(n586), .Z(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U655 ( .A1(G72), .A2(n616), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G85), .A2(n805), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G60), .A2(n634), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT66), .B(n591), .Z(n592) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n617), .A2(G47), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(G290) );
  NAND2_X1 U663 ( .A1(n706), .A2(G138), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G114), .A2(n901), .ZN(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT91), .B(n596), .Z(n602) );
  NAND2_X1 U666 ( .A1(G102), .A2(n909), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G126), .A2(n902), .ZN(n599) );
  AND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U670 ( .A(n705), .ZN(n605) );
  INV_X1 U671 ( .A(n685), .ZN(n607) );
  NOR2_X1 U672 ( .A1(G2084), .A2(n674), .ZN(n682) );
  NAND2_X1 U673 ( .A1(n607), .A2(n519), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n608), .B(KEYINPUT30), .ZN(n609) );
  NOR2_X1 U675 ( .A1(n609), .A2(G168), .ZN(n614) );
  NOR2_X1 U676 ( .A1(n657), .A2(G1961), .ZN(n610) );
  XOR2_X1 U677 ( .A(KEYINPUT93), .B(n610), .Z(n612) );
  XOR2_X1 U678 ( .A(G2078), .B(KEYINPUT25), .Z(n1009) );
  NOR2_X1 U679 ( .A1(n1009), .A2(n674), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n669) );
  AND2_X1 U681 ( .A1(G301), .A2(n669), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G79), .A2(n616), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G54), .A2(n617), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U686 ( .A(n620), .B(KEYINPUT76), .ZN(n624) );
  NAND2_X1 U687 ( .A1(G92), .A2(n805), .ZN(n622) );
  NAND2_X1 U688 ( .A1(G66), .A2(n634), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n626) );
  INV_X1 U691 ( .A(KEYINPUT15), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n626), .B(n625), .ZN(n627) );
  XOR2_X1 U693 ( .A(KEYINPUT77), .B(n627), .Z(n786) );
  INV_X1 U694 ( .A(n786), .ZN(n781) );
  NAND2_X1 U695 ( .A1(n805), .A2(G81), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G68), .A2(n616), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT13), .ZN(n633) );
  NAND2_X1 U700 ( .A1(G43), .A2(n617), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U702 ( .A1(G56), .A2(n634), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n635), .B(KEYINPUT14), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n636), .B(KEYINPUT75), .ZN(n637) );
  INV_X1 U705 ( .A(n937), .ZN(n801) );
  NOR2_X1 U706 ( .A1(n781), .A2(n801), .ZN(n644) );
  INV_X1 U707 ( .A(KEYINPUT96), .ZN(n643) );
  NAND2_X1 U708 ( .A1(G1996), .A2(n657), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT26), .ZN(n641) );
  NAND2_X1 U710 ( .A1(G1341), .A2(n674), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n650) );
  NAND2_X1 U713 ( .A1(n644), .A2(n650), .ZN(n649) );
  NAND2_X1 U714 ( .A1(G1348), .A2(n674), .ZN(n646) );
  NAND2_X1 U715 ( .A1(G2067), .A2(n657), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U717 ( .A(KEYINPUT97), .B(n647), .Z(n648) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n650), .A2(n937), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n651), .A2(n781), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n661) );
  INV_X1 U722 ( .A(G299), .ZN(n663) );
  NAND2_X1 U723 ( .A1(G2072), .A2(n657), .ZN(n656) );
  XOR2_X1 U724 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT94), .B(n654), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(n659) );
  INV_X1 U727 ( .A(G1956), .ZN(n864) );
  NOR2_X1 U728 ( .A1(n657), .A2(n864), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U733 ( .A(n664), .B(KEYINPUT28), .Z(n665) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT29), .ZN(n668) );
  INV_X1 U736 ( .A(n668), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n670), .A2(n518), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n517), .A2(n671), .ZN(n683) );
  NAND2_X1 U739 ( .A1(n683), .A2(G286), .ZN(n680) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n741), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT98), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G166), .A2(n673), .ZN(n677) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(KEYINPUT99), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U746 ( .A1(n606), .A2(n678), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(G8), .ZN(n687) );
  INV_X1 U749 ( .A(n683), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n735) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n698) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n698), .A2(n690), .ZN(n941) );
  NAND2_X1 U756 ( .A1(n735), .A2(n941), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n691), .B(KEYINPUT101), .ZN(n694) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n936) );
  INV_X1 U759 ( .A(n936), .ZN(n692) );
  OR2_X1 U760 ( .A1(n741), .A2(n692), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n695), .B(KEYINPUT64), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT102), .ZN(n701) );
  NAND2_X1 U765 ( .A1(n698), .A2(KEYINPUT33), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n741), .A2(n699), .ZN(n700) );
  NOR2_X2 U767 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n703), .B(n702), .ZN(n734) );
  XOR2_X1 U769 ( .A(G1981), .B(G305), .Z(n924) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n761) );
  XNOR2_X1 U771 ( .A(KEYINPUT37), .B(G2067), .ZN(n751) );
  BUF_X1 U772 ( .A(n706), .Z(n906) );
  NAND2_X1 U773 ( .A1(G140), .A2(n906), .ZN(n708) );
  NAND2_X1 U774 ( .A1(G104), .A2(n909), .ZN(n707) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(KEYINPUT34), .B(n709), .ZN(n715) );
  NAND2_X1 U777 ( .A1(G116), .A2(n901), .ZN(n711) );
  NAND2_X1 U778 ( .A1(G128), .A2(n902), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U780 ( .A(KEYINPUT92), .B(n712), .Z(n713) );
  XNOR2_X1 U781 ( .A(KEYINPUT35), .B(n713), .ZN(n714) );
  NOR2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U783 ( .A(KEYINPUT36), .B(n716), .ZN(n898) );
  NOR2_X1 U784 ( .A1(n751), .A2(n898), .ZN(n986) );
  NAND2_X1 U785 ( .A1(n761), .A2(n986), .ZN(n758) );
  NAND2_X1 U786 ( .A1(G141), .A2(n906), .ZN(n718) );
  NAND2_X1 U787 ( .A1(G129), .A2(n902), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n909), .A2(G105), .ZN(n719) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n719), .Z(n720) );
  NOR2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n901), .A2(G117), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n894) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n894), .ZN(n731) );
  NAND2_X1 U795 ( .A1(G131), .A2(n906), .ZN(n725) );
  NAND2_X1 U796 ( .A1(G119), .A2(n902), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G107), .A2(n901), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G95), .A2(n909), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n883) );
  NAND2_X1 U802 ( .A1(G1991), .A2(n883), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n982) );
  NAND2_X1 U804 ( .A1(n761), .A2(n982), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n758), .A2(n754), .ZN(n745) );
  INV_X1 U806 ( .A(n745), .ZN(n732) );
  AND2_X1 U807 ( .A1(n924), .A2(n732), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n747) );
  NOR2_X1 U809 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U810 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n735), .A2(n737), .ZN(n738) );
  AND2_X1 U812 ( .A1(n738), .A2(n741), .ZN(n743) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U814 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  NOR2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  OR2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n748), .B(KEYINPUT104), .ZN(n750) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n943) );
  NAND2_X1 U821 ( .A1(n943), .A2(n761), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n764) );
  NAND2_X1 U823 ( .A1(n751), .A2(n898), .ZN(n994) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n752) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n883), .ZN(n980) );
  NOR2_X1 U826 ( .A1(n752), .A2(n980), .ZN(n753) );
  XNOR2_X1 U827 ( .A(KEYINPUT105), .B(n753), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  OR2_X1 U829 ( .A1(n894), .A2(G1996), .ZN(n976) );
  NAND2_X1 U830 ( .A1(n756), .A2(n976), .ZN(n757) );
  XOR2_X1 U831 ( .A(KEYINPUT39), .B(n757), .Z(n759) );
  NAND2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n994), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U837 ( .A(G2438), .B(G2454), .Z(n767) );
  XNOR2_X1 U838 ( .A(G2435), .B(G2430), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U840 ( .A(n768), .B(G2427), .Z(n770) );
  XNOR2_X1 U841 ( .A(G1341), .B(G1348), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n770), .B(n769), .ZN(n774) );
  XOR2_X1 U843 ( .A(G2443), .B(G2446), .Z(n772) );
  XNOR2_X1 U844 ( .A(KEYINPUT106), .B(G2451), .ZN(n771) );
  XNOR2_X1 U845 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U846 ( .A(n774), .B(n773), .Z(n775) );
  AND2_X1 U847 ( .A1(G14), .A2(n775), .ZN(G401) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  BUF_X1 U849 ( .A(n776), .Z(G164) );
  NAND2_X1 U850 ( .A1(G94), .A2(G452), .ZN(n777) );
  XOR2_X1 U851 ( .A(KEYINPUT70), .B(n777), .Z(G173) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U853 ( .A(n778), .B(KEYINPUT74), .ZN(n779) );
  XOR2_X1 U854 ( .A(KEYINPUT10), .B(n779), .Z(n841) );
  NAND2_X1 U855 ( .A1(n841), .A2(G567), .ZN(n780) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n780), .Z(G234) );
  NAND2_X1 U857 ( .A1(n937), .A2(G860), .ZN(G153) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n783) );
  INV_X1 U859 ( .A(G868), .ZN(n822) );
  NAND2_X1 U860 ( .A1(n781), .A2(n822), .ZN(n782) );
  NAND2_X1 U861 ( .A1(n783), .A2(n782), .ZN(G284) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U863 ( .A1(G286), .A2(n822), .ZN(n784) );
  NOR2_X1 U864 ( .A1(n785), .A2(n784), .ZN(G297) );
  INV_X1 U865 ( .A(G860), .ZN(n803) );
  NAND2_X1 U866 ( .A1(n803), .A2(G559), .ZN(n787) );
  BUF_X1 U867 ( .A(n786), .Z(n928) );
  NAND2_X1 U868 ( .A1(n787), .A2(n928), .ZN(n788) );
  XNOR2_X1 U869 ( .A(n788), .B(KEYINPUT79), .ZN(n789) );
  XOR2_X1 U870 ( .A(KEYINPUT16), .B(n789), .Z(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n801), .ZN(n792) );
  NAND2_X1 U872 ( .A1(G868), .A2(n928), .ZN(n790) );
  NOR2_X1 U873 ( .A1(G559), .A2(n790), .ZN(n791) );
  NOR2_X1 U874 ( .A1(n792), .A2(n791), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n902), .ZN(n793) );
  XNOR2_X1 U876 ( .A(n793), .B(KEYINPUT18), .ZN(n795) );
  NAND2_X1 U877 ( .A1(n901), .A2(G111), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G135), .A2(n906), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G99), .A2(n909), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U882 ( .A1(n799), .A2(n798), .ZN(n979) );
  XNOR2_X1 U883 ( .A(G2096), .B(n979), .ZN(n800) );
  INV_X1 U884 ( .A(G2100), .ZN(n857) );
  NAND2_X1 U885 ( .A1(n800), .A2(n857), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G559), .A2(n928), .ZN(n802) );
  XOR2_X1 U887 ( .A(n802), .B(n801), .Z(n820) );
  NAND2_X1 U888 ( .A1(n803), .A2(n820), .ZN(n813) );
  NAND2_X1 U889 ( .A1(G67), .A2(n634), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n804), .B(KEYINPUT80), .ZN(n812) );
  NAND2_X1 U891 ( .A1(G80), .A2(n616), .ZN(n807) );
  NAND2_X1 U892 ( .A1(G93), .A2(n805), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U894 ( .A1(G55), .A2(n617), .ZN(n808) );
  XNOR2_X1 U895 ( .A(KEYINPUT81), .B(n808), .ZN(n809) );
  NOR2_X1 U896 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n812), .A2(n811), .ZN(n823) );
  XNOR2_X1 U898 ( .A(n813), .B(n823), .ZN(G145) );
  XOR2_X1 U899 ( .A(KEYINPUT87), .B(G166), .Z(n814) );
  XNOR2_X1 U900 ( .A(n814), .B(n823), .ZN(n817) );
  XOR2_X1 U901 ( .A(G299), .B(G290), .Z(n815) );
  XNOR2_X1 U902 ( .A(n815), .B(G288), .ZN(n816) );
  XNOR2_X1 U903 ( .A(n817), .B(n816), .ZN(n819) );
  XNOR2_X1 U904 ( .A(G305), .B(KEYINPUT19), .ZN(n818) );
  XNOR2_X1 U905 ( .A(n819), .B(n818), .ZN(n849) );
  XNOR2_X1 U906 ( .A(n820), .B(n849), .ZN(n821) );
  NAND2_X1 U907 ( .A1(n821), .A2(G868), .ZN(n825) );
  NAND2_X1 U908 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n827), .ZN(n828) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U914 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n831) );
  NAND2_X1 U917 ( .A1(G132), .A2(G82), .ZN(n830) );
  XNOR2_X1 U918 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U919 ( .A(n832), .B(KEYINPUT88), .ZN(n833) );
  NOR2_X1 U920 ( .A1(G218), .A2(n833), .ZN(n834) );
  NAND2_X1 U921 ( .A1(G96), .A2(n834), .ZN(n845) );
  NAND2_X1 U922 ( .A1(n845), .A2(G2106), .ZN(n838) );
  NAND2_X1 U923 ( .A1(G69), .A2(G120), .ZN(n835) );
  NOR2_X1 U924 ( .A1(G237), .A2(n835), .ZN(n836) );
  NAND2_X1 U925 ( .A1(G108), .A2(n836), .ZN(n846) );
  NAND2_X1 U926 ( .A1(n846), .A2(G567), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n838), .A2(n837), .ZN(n922) );
  NAND2_X1 U928 ( .A1(G661), .A2(G483), .ZN(n839) );
  XNOR2_X1 U929 ( .A(KEYINPUT90), .B(n839), .ZN(n840) );
  NOR2_X1 U930 ( .A1(n922), .A2(n840), .ZN(n844) );
  NAND2_X1 U931 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n841), .ZN(G217) );
  INV_X1 U933 ( .A(n841), .ZN(G223) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U935 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(G188) );
  NOR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(G325) );
  XNOR2_X1 U939 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U941 ( .A(G132), .ZN(G219) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G82), .ZN(G220) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  XOR2_X1 U946 ( .A(n928), .B(n937), .Z(n848) );
  XOR2_X1 U947 ( .A(G286), .B(G301), .Z(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  NOR2_X1 U950 ( .A1(G37), .A2(n851), .ZN(G397) );
  XOR2_X1 U951 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT108), .B(G2096), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n854), .B(KEYINPUT109), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2072), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n857), .B(G2084), .ZN(n859) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2090), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2678), .B(KEYINPUT43), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(G227) );
  XNOR2_X1 U963 ( .A(G1976), .B(n864), .ZN(n866) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1971), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(n867), .B(KEYINPUT41), .Z(n869) );
  XNOR2_X1 U967 ( .A(G1966), .B(G1981), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U969 ( .A(G2474), .B(G1961), .Z(n871) );
  XNOR2_X1 U970 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n902), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT44), .B(n874), .Z(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT111), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G112), .A2(n901), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G136), .A2(n906), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G100), .A2(n909), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(G162) );
  XOR2_X1 U982 ( .A(G164), .B(n979), .Z(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n884), .B(KEYINPUT113), .Z(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n897) );
  NAND2_X1 U987 ( .A1(G118), .A2(n901), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G130), .A2(n902), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G142), .A2(n906), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G106), .A2(n909), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(n891), .B(KEYINPUT45), .Z(n892) );
  NOR2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n898), .B(G162), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n914) );
  NAND2_X1 U999 ( .A1(G115), .A2(n901), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G127), .A2(n902), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(KEYINPUT47), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n906), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(n909), .A2(G103), .ZN(n910) );
  XOR2_X1 U1006 ( .A(KEYINPUT112), .B(n910), .Z(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n990) );
  XOR2_X1 U1008 ( .A(n990), .B(G160), .Z(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n917), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(G401), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT114), .B(n918), .Z(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n919), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n922), .ZN(G319) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1021 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n1029) );
  XNOR2_X1 U1022 ( .A(KEYINPUT56), .B(G16), .ZN(n947) );
  XNOR2_X1 U1023 ( .A(G168), .B(G1966), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT120), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT57), .ZN(n932) );
  XOR2_X1 U1027 ( .A(G299), .B(G1956), .Z(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT121), .ZN(n930) );
  XOR2_X1 U1029 ( .A(G1348), .B(n928), .Z(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n934) );
  XOR2_X1 U1032 ( .A(G1961), .B(G171), .Z(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n945) );
  NAND2_X1 U1034 ( .A1(G1971), .A2(G303), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1036 ( .A(G1341), .B(n937), .Z(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n973) );
  XNOR2_X1 U1042 ( .A(G1961), .B(G5), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n960) );
  XOR2_X1 U1045 ( .A(KEYINPUT122), .B(G4), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G1348), .B(KEYINPUT59), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n951), .B(n950), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G20), .B(G1956), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G6), .B(G1981), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT60), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT61), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT123), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(G16), .A2(n970), .ZN(n971) );
  XOR2_X1 U1066 ( .A(KEYINPUT124), .B(n971), .Z(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(KEYINPUT125), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(G11), .ZN(n1003) );
  XNOR2_X1 U1070 ( .A(G2090), .B(G162), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT51), .ZN(n988) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G160), .B(G2084), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n997) );
  XNOR2_X1 U1079 ( .A(G164), .B(G2078), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT115), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G2072), .B(n990), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT50), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1086 ( .A(KEYINPUT52), .B(n998), .Z(n999) );
  NOR2_X1 U1087 ( .A1(KEYINPUT55), .A2(n999), .ZN(n1000) );
  INV_X1 U1088 ( .A(G29), .ZN(n1004) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n1004), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT116), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1027) );
  XOR2_X1 U1092 ( .A(n1004), .B(KEYINPUT119), .Z(n1025) );
  XOR2_X1 U1093 ( .A(G2090), .B(G35), .Z(n1019) );
  XOR2_X1 U1094 ( .A(G2072), .B(G33), .Z(n1005) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(G28), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G25), .B(G1991), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT117), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G2067), .B(G26), .Z(n1008) );
  XOR2_X1 U1099 ( .A(G1996), .B(G32), .Z(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(G27), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT118), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT53), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G34), .B(G2084), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT54), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(KEYINPUT55), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(n1029), .B(n1028), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

