//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  NAND2_X1  g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT98), .B1(G71gat), .B2(G78gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n206), .A2(new_n203), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G71gat), .ZN(new_n210));
  INV_X1    g009(.A(G78gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n210), .B(new_n211), .C1(KEYINPUT99), .C2(KEYINPUT9), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n203), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n205), .A2(KEYINPUT99), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n202), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G231gat), .A2(G233gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT94), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G8gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  AOI21_X1  g025(.A(G1gat), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT95), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(KEYINPUT95), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(new_n217), .B2(new_n216), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n222), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G155gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(G183gat), .B(G211gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT7), .ZN(new_n243));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244));
  INV_X1    g043(.A(G85gat), .ZN(new_n245));
  INV_X1    g044(.A(G92gat), .ZN(new_n246));
  AOI22_X1  g045(.A1(KEYINPUT8), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G99gat), .B(G106gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT100), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n243), .A2(KEYINPUT100), .A3(new_n249), .A4(new_n247), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT15), .ZN(new_n258));
  NOR3_X1   g057(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT92), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(G29gat), .B2(G36gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G29gat), .A2(G36gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n261), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT15), .A3(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n254), .A2(new_n268), .B1(KEYINPUT41), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(KEYINPUT93), .B(KEYINPUT17), .C1(new_n263), .C2(new_n267), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n254), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n272), .B2(new_n268), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n270), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G190gat), .B(G218gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT101), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n269), .A2(KEYINPUT41), .ZN(new_n282));
  XNOR2_X1  g081(.A(G134gat), .B(G162gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n280), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n285), .B(new_n270), .C1(new_n275), .C2(new_n277), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n281), .B2(new_n286), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n241), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n292));
  INV_X1    g091(.A(new_n216), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n252), .B2(new_n253), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n250), .A2(new_n216), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n254), .A2(KEYINPUT10), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT102), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(KEYINPUT102), .A3(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n294), .A2(new_n301), .A3(new_n295), .ZN(new_n304));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n301), .B(KEYINPUT103), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n296), .B2(new_n297), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n312), .B2(new_n304), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n291), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n317));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n268), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n230), .B2(new_n231), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n228), .A2(KEYINPUT95), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n268), .A3(new_n229), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n228), .B1(new_n320), .B2(KEYINPUT17), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n274), .B2(new_n273), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n318), .A3(new_n323), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT18), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G197gat), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT11), .B(G169gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n327), .A2(new_n328), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n329), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G15gat), .B(G43gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G227gat), .ZN(new_n344));
  INV_X1    g143(.A(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  INV_X1    g147(.A(G183gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT68), .B1(new_n349), .B2(KEYINPUT27), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(G183gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n352), .B2(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n348), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n362), .B(new_n348), .C1(new_n355), .C2(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(KEYINPUT27), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n352), .A2(G183gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT28), .A4(new_n358), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(KEYINPUT26), .ZN(new_n369));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n368), .B2(KEYINPUT26), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n369), .A2(new_n372), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n368), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT25), .B1(new_n374), .B2(KEYINPUT23), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n368), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n379), .B(new_n370), .C1(new_n368), .C2(new_n376), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n349), .A2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n358), .A2(G183gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(G183gat), .A3(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT66), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT66), .ZN(new_n389));
  XNOR2_X1  g188(.A(G183gat), .B(G190gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n389), .B(new_n386), .C1(new_n390), .C2(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(new_n384), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT24), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n371), .B1(new_n368), .B2(new_n376), .ZN(new_n396));
  OR2_X1    g195(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(G169gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n397), .A2(KEYINPUT23), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(new_n396), .A3(new_n386), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n367), .A2(new_n373), .B1(new_n393), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G120gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G113gat), .ZN(new_n408));
  INV_X1    g207(.A(G113gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G120gat), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT1), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI211_X1 g212(.A(KEYINPUT71), .B(KEYINPUT1), .C1(new_n408), .C2(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT71), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(new_n405), .C1(new_n412), .C2(new_n411), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(new_n373), .ZN(new_n422));
  INV_X1    g221(.A(new_n366), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n360), .B2(KEYINPUT69), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n424), .B2(new_n363), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n381), .A2(new_n392), .B1(new_n402), .B2(new_n401), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n347), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n343), .B1(new_n428), .B2(KEYINPUT33), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(KEYINPUT32), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n420), .A2(new_n347), .A3(new_n427), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(KEYINPUT34), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(KEYINPUT32), .A3(new_n430), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n438), .B2(new_n431), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  OAI22_X1  g241(.A1(new_n438), .A2(new_n431), .B1(new_n442), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n437), .B2(new_n442), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n367), .A2(new_n373), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n393), .A2(new_n403), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n425), .B2(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(G226gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT29), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456));
  INV_X1    g255(.A(G211gat), .ZN(new_n457));
  INV_X1    g256(.A(G218gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(KEYINPUT22), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G211gat), .B(G218gat), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n460), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n404), .A2(new_n453), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n455), .A2(KEYINPUT74), .A3(new_n463), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT75), .B(new_n452), .C1(new_n404), .C2(KEYINPUT29), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n460), .B(new_n461), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT29), .B1(new_n447), .B2(new_n448), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n453), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n474), .A3(new_n470), .A4(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT76), .ZN(new_n480));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n481), .B(new_n482), .Z(new_n483));
  NAND4_X1  g282(.A1(new_n469), .A2(new_n478), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT77), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n478), .A3(new_n480), .ZN(new_n491));
  INV_X1    g290(.A(new_n483), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n485), .B2(new_n484), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(G141gat), .ZN(new_n501));
  INV_X1    g300(.A(G148gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G141gat), .A2(G148gat), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G162gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G155gat), .ZN(new_n507));
  INV_X1    g306(.A(G155gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G162gat), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT2), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n505), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n503), .A2(new_n514), .A3(new_n504), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(new_n509), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n516), .A2(KEYINPUT78), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT78), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT3), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(KEYINPUT78), .A3(new_n517), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n515), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n528), .A3(new_n421), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT80), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n520), .A2(KEYINPUT3), .B1(new_n415), .B2(new_n418), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT80), .B1(new_n532), .B2(new_n528), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n500), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n421), .B2(new_n520), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT79), .B(G155gat), .Z(new_n538));
  OAI21_X1  g337(.A(KEYINPUT2), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  AND4_X1   g338(.A1(new_n503), .A2(new_n507), .A3(new_n509), .A4(new_n504), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n524), .A2(new_n525), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n541), .A2(new_n418), .A3(new_n415), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n499), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n500), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n530), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n532), .A2(KEYINPUT80), .A3(new_n528), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n545), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n421), .A2(new_n520), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n418), .A3(new_n415), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n500), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT83), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT5), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n421), .A2(new_n520), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n418), .A2(new_n415), .B1(new_n526), .B2(new_n515), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n547), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT83), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n535), .A3(new_n418), .A4(new_n415), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT82), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n419), .A2(new_n565), .A3(new_n535), .A4(new_n541), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n554), .A2(new_n543), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n546), .A2(new_n552), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G1gat), .B(G29gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT0), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G85gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  AOI21_X1  g373(.A(new_n498), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n570), .A2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n497), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n546), .A2(new_n552), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n555), .A2(new_n556), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n537), .B1(new_n560), .B2(KEYINPUT83), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n579), .B(new_n580), .C1(new_n534), .C2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(new_n498), .A3(new_n574), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n497), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n534), .A2(new_n499), .A3(new_n545), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT84), .B1(new_n550), .B2(new_n551), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n574), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n577), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n496), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT29), .B1(new_n541), .B2(new_n527), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n474), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT3), .B1(new_n474), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n541), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT86), .B1(new_n596), .B2(new_n541), .ZN(new_n599));
  NAND2_X1  g398(.A1(G228gat), .A2(G233gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n600), .B(new_n599), .C1(new_n594), .C2(new_n597), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G22gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G78gat), .B(G106gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT31), .B(G50gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n604), .A2(new_n605), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT87), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  INV_X1    g412(.A(new_n610), .ZN(new_n614));
  OAI21_X1  g413(.A(G22gat), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n611), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n446), .B1(new_n592), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n455), .A2(new_n474), .A3(new_n464), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(KEYINPUT37), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n472), .A2(new_n463), .A3(new_n477), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT38), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(new_n492), .C1(new_n491), .C2(KEYINPUT37), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n582), .B(new_n574), .C1(new_n585), .C2(new_n586), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT6), .B1(new_n627), .B2(new_n589), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n583), .A2(new_n497), .B1(new_n588), .B2(new_n587), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n484), .B(new_n625), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n492), .A2(KEYINPUT37), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n493), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n491), .A2(KEYINPUT37), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n618), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n536), .A2(new_n544), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n548), .B2(new_n549), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n500), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n588), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n558), .A2(new_n559), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n643), .B2(new_n500), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(new_n639), .B2(new_n500), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n576), .B1(new_n637), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(KEYINPUT40), .A3(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT88), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT88), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n642), .A2(new_n650), .A3(KEYINPUT40), .A4(new_n645), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n490), .B2(new_n495), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n620), .B1(new_n636), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n484), .A2(new_n488), .A3(new_n485), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n488), .B1(new_n484), .B2(new_n485), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n652), .B(new_n647), .C1(new_n658), .C2(new_n494), .ZN(new_n659));
  INV_X1    g458(.A(new_n634), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n492), .B1(new_n491), .B2(KEYINPUT37), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT38), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(new_n591), .A3(new_n484), .A4(new_n625), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n659), .A2(new_n663), .A3(KEYINPUT89), .A4(new_n618), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n619), .B1(new_n655), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n658), .A2(new_n494), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT35), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n618), .A2(new_n440), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n591), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT90), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n592), .A2(KEYINPUT90), .A3(new_n668), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n444), .A2(new_n618), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n592), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n672), .A2(new_n673), .B1(new_n675), .B2(KEYINPUT35), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n340), .B1(new_n665), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(KEYINPUT35), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n655), .A2(new_n664), .ZN(new_n682));
  INV_X1    g481(.A(new_n446), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n669), .ZN(new_n684));
  INV_X1    g483(.A(new_n618), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT97), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n340), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n316), .B1(new_n678), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n591), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  INV_X1    g492(.A(new_n691), .ZN(new_n694));
  INV_X1    g493(.A(G8gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n226), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n697));
  NOR4_X1   g496(.A1(new_n694), .A2(new_n666), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n691), .B2(new_n496), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(KEYINPUT42), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g500(.A(new_n440), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n694), .A2(G15gat), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n694), .B2(new_n446), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n691), .A2(new_n685), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NOR2_X1   g507(.A1(new_n240), .A2(new_n314), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n339), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n289), .A2(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n687), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT104), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(new_n681), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n289), .B1(new_n681), .B2(new_n687), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n591), .B(new_n711), .C1(new_n718), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n676), .B1(new_n715), .B2(new_n716), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n725), .A2(new_n713), .B1(new_n720), .B2(new_n719), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n591), .A4(new_n711), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(G29gat), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n678), .A2(new_n690), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n289), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G29gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n591), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT45), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n730), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n678), .B2(new_n690), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(new_n737), .A3(new_n732), .A4(new_n591), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n728), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1328gat));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n666), .A2(G36gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n736), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n736), .A2(new_n750), .A3(new_n746), .A4(new_n747), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n726), .A2(new_n711), .ZN(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n753), .B2(new_n666), .ZN(new_n754));
  INV_X1    g553(.A(new_n747), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT46), .B1(new_n731), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n745), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n749), .A2(new_n751), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(KEYINPUT108), .A3(new_n754), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1329gat));
  NAND3_X1  g560(.A1(new_n726), .A2(new_n683), .A3(new_n711), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n702), .A2(G43gat), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n736), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(KEYINPUT109), .B(KEYINPUT47), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n762), .A2(G43gat), .B1(new_n736), .B2(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n766), .A2(new_n770), .ZN(G1330gat));
  AOI21_X1  g570(.A(new_n618), .B1(new_n736), .B2(KEYINPUT110), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n731), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(G50gat), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n753), .A2(new_n776), .A3(new_n618), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT48), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT48), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1331gat));
  NAND2_X1  g579(.A1(new_n717), .A2(new_n681), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n340), .A2(new_n241), .A3(new_n290), .A4(new_n315), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n591), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g585(.A1(new_n783), .A2(new_n666), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  OR3_X1    g590(.A1(new_n783), .A2(KEYINPUT111), .A3(new_n702), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT111), .B1(new_n783), .B2(new_n702), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n210), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n784), .A2(G71gat), .A3(new_n683), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1334gat));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n618), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(new_n211), .ZN(G1335gat));
  NOR3_X1   g601(.A1(new_n340), .A2(new_n240), .A3(new_n289), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n781), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n245), .A3(new_n591), .A4(new_n314), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n340), .A2(new_n240), .A3(new_n315), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n726), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n591), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n245), .ZN(G1336gat));
  NOR3_X1   g611(.A1(new_n666), .A2(G92gat), .A3(new_n315), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n246), .B1(new_n810), .B2(new_n496), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n807), .A2(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n810), .A2(new_n496), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n246), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1337gat));
  INV_X1    g620(.A(G99gat), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n822), .A3(new_n440), .A4(new_n314), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n810), .A2(new_n683), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n822), .ZN(G1338gat));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n685), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n618), .A2(G106gat), .A3(new_n315), .ZN(new_n828));
  INV_X1    g627(.A(new_n806), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n804), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n827), .A2(KEYINPUT112), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n831), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n834));
  INV_X1    g633(.A(G106gat), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n810), .B2(new_n685), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n837), .ZN(G1339gat));
  NAND3_X1  g637(.A1(new_n291), .A2(new_n339), .A3(new_n315), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n296), .A2(new_n297), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n311), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n303), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n307), .B1(new_n312), .B2(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT55), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n310), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n321), .A2(new_n323), .A3(new_n319), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n318), .B1(new_n326), .B2(new_n323), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n333), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n850), .B(new_n853), .C1(new_n287), .C2(new_n288), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n314), .A3(new_n853), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n849), .B2(new_n339), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n857), .B2(new_n289), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n839), .B1(new_n858), .B2(new_n240), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n591), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n666), .A2(new_n674), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT114), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n409), .A3(new_n340), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n685), .A2(new_n702), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n496), .A2(new_n669), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n339), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(G1340gat));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n407), .A3(new_n314), .ZN(new_n870));
  OAI21_X1  g669(.A(G120gat), .B1(new_n867), .B2(new_n315), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1341gat));
  OR3_X1    g671(.A1(new_n867), .A2(new_n221), .A3(new_n241), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n221), .B1(new_n862), .B2(new_n241), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(KEYINPUT115), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G1342gat));
  OR3_X1    g676(.A1(new_n862), .A2(G134gat), .A3(new_n289), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n867), .B2(new_n289), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n683), .A2(new_n618), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n860), .A2(new_n666), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n501), .A3(new_n340), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n859), .A2(new_n886), .A3(new_n685), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n446), .A3(new_n866), .ZN(new_n888));
  INV_X1    g687(.A(new_n855), .ZN(new_n889));
  INV_X1    g688(.A(new_n856), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n848), .A2(new_n310), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n312), .A2(new_n840), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n308), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n303), .B2(new_n842), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n895), .B2(KEYINPUT55), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n845), .A2(KEYINPUT116), .A3(new_n846), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n339), .B1(new_n898), .B2(KEYINPUT117), .ZN(new_n899));
  INV_X1    g698(.A(new_n891), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n895), .A2(new_n892), .A3(KEYINPUT55), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT116), .B1(new_n845), .B2(new_n846), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n890), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n889), .B1(new_n906), .B2(new_n290), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n241), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n839), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n685), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n888), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n340), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n885), .B1(new_n912), .B2(new_n501), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n884), .A2(new_n502), .A3(new_n314), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n866), .A2(new_n446), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n315), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n839), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n907), .B2(new_n241), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n886), .B1(new_n921), .B2(new_n618), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n859), .A2(KEYINPUT57), .A3(new_n685), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n922), .A2(KEYINPUT119), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n909), .B2(new_n685), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n502), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n924), .A2(new_n925), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n927), .B2(new_n928), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n922), .A2(KEYINPUT119), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n918), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT120), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n916), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT59), .B(new_n502), .C1(new_n911), .C2(new_n314), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n915), .B1(new_n938), .B2(new_n939), .ZN(G1345gat));
  NOR2_X1   g739(.A1(new_n241), .A2(new_n538), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n884), .A2(new_n240), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n911), .A2(new_n941), .B1(new_n538), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT121), .Z(G1346gat));
  AOI21_X1  g743(.A(G162gat), .B1(new_n884), .B2(new_n290), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n289), .A2(new_n506), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n911), .B2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n666), .A2(new_n591), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n859), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(new_n674), .ZN(new_n950));
  AOI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n340), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n865), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n339), .A2(new_n398), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G1348gat));
  AOI21_X1  g755(.A(G176gat), .B1(new_n950), .B2(new_n314), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n315), .B1(new_n397), .B2(new_n399), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n954), .B2(new_n958), .ZN(G1349gat));
  NAND2_X1  g758(.A1(new_n954), .A2(new_n240), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT123), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n954), .A2(new_n962), .A3(new_n240), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(G183gat), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n950), .A2(new_n364), .A3(new_n365), .A4(new_n240), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT60), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1350gat));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n290), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT61), .B1(new_n971), .B2(G190gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n358), .A3(new_n290), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT124), .ZN(new_n975));
  OR3_X1    g774(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n949), .A2(new_n883), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT125), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n340), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n926), .A2(new_n929), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n683), .A2(new_n591), .A3(new_n666), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n340), .A2(G197gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G1352gat));
  OAI21_X1  g784(.A(G204gat), .B1(new_n982), .B2(new_n315), .ZN(new_n986));
  AOI21_X1  g785(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n949), .A2(new_n314), .A3(new_n883), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n978), .A2(new_n457), .A3(new_n240), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n980), .A2(new_n240), .A3(new_n981), .ZN(new_n994));
  AND4_X1   g793(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT63), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n457), .B1(KEYINPUT127), .B2(new_n996), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n994), .A2(new_n997), .B1(new_n993), .B2(KEYINPUT63), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n992), .B1(new_n995), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n982), .B2(new_n289), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n978), .A2(new_n458), .A3(new_n290), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


