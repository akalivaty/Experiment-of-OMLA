//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n203), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XNOR2_X1  g0021(.A(G238), .B(G244), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT2), .B(G226), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n225), .B(new_n228), .ZN(G358));
  XOR2_X1   g0029(.A(G87), .B(G97), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G107), .B(G116), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G68), .B(G77), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G351));
  NAND3_X1  g0038(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n239));
  INV_X1    g0039(.A(KEYINPUT68), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n239), .A2(new_n240), .A3(new_n209), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g0042(.A(new_n240), .B1(new_n239), .B2(new_n209), .ZN(new_n243));
  INV_X1    g0043(.A(G13), .ZN(new_n244));
  NOR3_X1   g0044(.A1(new_n244), .A2(new_n210), .A3(G1), .ZN(new_n245));
  NOR3_X1   g0045(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT15), .B(G87), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n246), .A2(KEYINPUT86), .A3(new_n248), .A4(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT86), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n239), .A2(new_n209), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n244), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(new_n241), .A4(new_n251), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n258), .B2(new_n247), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n210), .B(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT85), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT85), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(new_n210), .A4(G68), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G97), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT19), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n210), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G97), .A2(G107), .ZN(new_n274));
  INV_X1    g0074(.A(G87), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G97), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(new_n249), .B2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n210), .A2(KEYINPUT69), .A3(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(KEYINPUT19), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n254), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n247), .A2(new_n245), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n260), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT87), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n264), .A2(new_n269), .ZN(new_n288));
  INV_X1    g0088(.A(new_n281), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT69), .B1(new_n210), .B2(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(G97), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n272), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n277), .A3(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(new_n254), .B1(new_n245), .B2(new_n247), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT87), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(new_n260), .ZN(new_n296));
  OAI211_X1 g0096(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(G238), .B(new_n298), .C1(new_n261), .C2(new_n262), .ZN(new_n299));
  INV_X1    g0099(.A(G116), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n297), .B(new_n299), .C1(new_n249), .C2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n209), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT66), .B1(new_n302), .B2(new_n209), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT66), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(G1), .A4(G13), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G45), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT83), .B1(new_n310), .B2(G1), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT83), .ZN(new_n312));
  INV_X1    g0112(.A(G1), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(G45), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n314), .A3(G250), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT84), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n310), .A2(G1), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n305), .A2(G274), .A3(new_n308), .A4(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n311), .A2(new_n314), .A3(G250), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT84), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n305), .A4(new_n308), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n304), .A2(new_n316), .A3(new_n318), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n316), .A2(new_n321), .A3(new_n318), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n304), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n287), .A2(new_n296), .A3(new_n324), .A4(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT88), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n246), .A2(new_n329), .A3(G87), .A4(new_n251), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT88), .B1(new_n258), .B2(new_n275), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n284), .A3(new_n285), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n322), .A2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G1698), .B1(new_n265), .B2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G222), .ZN(new_n341));
  INV_X1    g0141(.A(G77), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n267), .A2(G1698), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n341), .B1(new_n342), .B2(new_n267), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n305), .A2(G274), .A3(new_n308), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n313), .B1(G41), .B2(G45), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n345), .A2(new_n303), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n305), .A2(new_n308), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT67), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n305), .A2(new_n352), .A3(new_n308), .A4(new_n347), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G226), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n255), .A2(new_n241), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n289), .A2(new_n290), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT8), .B(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G20), .A2(G33), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n365), .A2(new_n367), .B1(new_n368), .B2(new_n210), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n361), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n313), .A2(G20), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n246), .A2(G50), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G50), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n245), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n370), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n357), .B1(new_n334), .B2(new_n356), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n360), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n378), .B(KEYINPUT9), .ZN(new_n383));
  INV_X1    g0183(.A(new_n381), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n359), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n305), .A2(new_n348), .A3(G274), .A4(new_n308), .ZN(new_n387));
  INV_X1    g0187(.A(G238), .ZN(new_n388));
  INV_X1    g0188(.A(G107), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n344), .A2(new_n388), .B1(new_n389), .B2(new_n267), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n340), .A2(new_n391), .A3(G232), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n340), .A2(G232), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT71), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n303), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n387), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n354), .A2(G244), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n323), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n362), .A2(new_n247), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n363), .A2(new_n367), .B1(new_n210), .B2(new_n342), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n254), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G77), .B2(new_n257), .ZN(new_n404));
  INV_X1    g0204(.A(new_n254), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT72), .B1(new_n405), .B2(new_n257), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT72), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n245), .A2(new_n254), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n371), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n342), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n394), .A2(new_n392), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n303), .B1(new_n413), .B2(new_n390), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(new_n326), .A3(new_n387), .A4(new_n398), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n400), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G200), .B1(new_n397), .B2(new_n399), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(G190), .A3(new_n387), .A4(new_n398), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n356), .A2(new_n323), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n349), .A2(new_n326), .A3(new_n355), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n378), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n386), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT75), .B(KEYINPUT14), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n354), .A2(G238), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G226), .A2(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G232), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(G1698), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n267), .B1(G33), .B2(G97), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n387), .B1(new_n431), .B2(new_n396), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n426), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n388), .B1(new_n351), .B2(new_n353), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n435), .A2(KEYINPUT13), .A3(new_n432), .ZN(new_n436));
  OAI211_X1 g0236(.A(G169), .B(new_n425), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n427), .A2(new_n426), .A3(new_n433), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT13), .B1(new_n435), .B2(new_n432), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n323), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT74), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n434), .B2(new_n436), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT14), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n441), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n362), .A2(new_n342), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n367), .A2(new_n373), .B1(new_n210), .B2(G68), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n361), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT11), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G68), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n409), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n245), .A2(new_n454), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n448), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n438), .A2(new_n439), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G200), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n460), .B(new_n464), .C1(new_n334), .C2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n363), .B1(new_n313), .B2(G20), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n246), .A2(new_n468), .B1(new_n245), .B2(new_n363), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n261), .A2(new_n262), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT7), .B1(new_n471), .B2(new_n210), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT7), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n261), .A2(new_n262), .A3(new_n473), .A4(G20), .ZN(new_n474));
  OAI21_X1  g0274(.A(G68), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(G58), .B(G68), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(G20), .B1(G159), .B2(new_n366), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT16), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n405), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT76), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n265), .A2(new_n481), .A3(new_n266), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT76), .B1(new_n261), .B2(new_n262), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n210), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n474), .B1(new_n484), .B2(new_n473), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT16), .B(new_n477), .C1(new_n485), .C2(new_n454), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n470), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n387), .B1(new_n350), .B2(new_n429), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT80), .A2(G190), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT80), .A2(G190), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G87), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT77), .ZN(new_n495));
  OAI211_X1 g0295(.A(G223), .B(new_n298), .C1(new_n261), .C2(new_n262), .ZN(new_n496));
  OAI211_X1 g0296(.A(G226), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n303), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT78), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n387), .B(new_n500), .C1(new_n350), .C2(new_n429), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n489), .A2(new_n493), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G200), .ZN(new_n503));
  INV_X1    g0303(.A(new_n499), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n488), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n487), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT17), .B1(new_n487), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n467), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n487), .A2(new_n506), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n487), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(KEYINPUT81), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT18), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n489), .A2(new_n326), .A3(new_n499), .A4(new_n501), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n323), .B1(new_n504), .B2(new_n488), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n487), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n487), .A2(new_n518), .A3(new_n515), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(KEYINPUT79), .ZN(new_n521));
  INV_X1    g0321(.A(new_n487), .ZN(new_n522));
  INV_X1    g0322(.A(new_n518), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT79), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n509), .A2(new_n514), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n424), .A2(new_n466), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n389), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(G97), .B(G107), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n534), .A2(new_n210), .B1(new_n342), .B2(new_n367), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n473), .B1(new_n267), .B2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n471), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n389), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n254), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n258), .A2(new_n278), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n257), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n298), .C1(new_n261), .C2(new_n262), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT4), .B1(new_n340), .B2(G244), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n303), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  INV_X1    g0352(.A(G41), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT5), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT5), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT82), .B1(new_n555), .B2(G41), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(G41), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n317), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n346), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n558), .A2(G257), .A3(new_n305), .A4(new_n308), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n551), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n326), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n305), .A2(G274), .A3(new_n308), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n559), .A2(new_n309), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(G257), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n323), .B1(new_n567), .B2(new_n551), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n544), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n472), .B2(new_n474), .ZN(new_n570));
  AND2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n533), .B1(new_n571), .B2(new_n274), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n530), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n366), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n405), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n575), .A2(new_n540), .A3(new_n542), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n562), .A2(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n567), .A2(G190), .A3(new_n551), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n569), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n210), .A2(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT91), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n256), .B(new_n581), .C1(new_n582), .C2(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(KEYINPUT25), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n389), .B2(new_n258), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n210), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n267), .A2(new_n589), .A3(new_n210), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n249), .A2(new_n300), .A3(G20), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT89), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT23), .B1(new_n581), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI211_X1 g0396(.A(KEYINPUT89), .B(new_n596), .C1(new_n210), .C2(G107), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n591), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n591), .B2(new_n598), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n254), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT90), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n591), .A2(new_n592), .A3(new_n598), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n254), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n586), .B1(new_n602), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(new_n298), .C1(new_n261), .C2(new_n262), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G33), .A2(G294), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n303), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n558), .A2(G264), .A3(new_n305), .A4(new_n308), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n560), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n503), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT93), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT92), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n618), .B2(G190), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n616), .A2(new_n617), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT92), .A3(new_n334), .A4(new_n560), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n621), .A2(new_n623), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n580), .B1(new_n611), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n250), .A2(new_n300), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n406), .B2(new_n408), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n256), .A2(G20), .A3(new_n300), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n545), .B(new_n210), .C1(G33), .C2(new_n278), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n300), .A2(G20), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n254), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n632), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n640));
  OAI211_X1 g0440(.A(G257), .B(new_n298), .C1(new_n261), .C2(new_n262), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n303), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n558), .A2(G270), .A3(new_n305), .A4(new_n308), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n560), .A2(new_n644), .A3(new_n645), .A4(new_n492), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n560), .A2(new_n644), .A3(new_n645), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n639), .B(new_n646), .C1(new_n648), .C2(new_n503), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n630), .A2(new_n638), .A3(new_n631), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(G169), .A3(new_n647), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT21), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(G179), .A3(new_n650), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n650), .A2(new_n647), .A3(KEYINPUT21), .A4(G169), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n649), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n586), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n609), .B1(new_n608), .B2(new_n254), .ZN(new_n658));
  AOI211_X1 g0458(.A(KEYINPUT90), .B(new_n405), .C1(new_n606), .C2(new_n607), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n618), .A2(G179), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n323), .B2(new_n618), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n656), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n339), .A2(new_n529), .A3(new_n628), .A4(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n423), .ZN(new_n665));
  INV_X1    g0465(.A(new_n520), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n519), .ZN(new_n667));
  INV_X1    g0467(.A(new_n416), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n461), .B1(new_n465), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n509), .A2(new_n514), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n672), .B2(new_n386), .ZN(new_n673));
  INV_X1    g0473(.A(new_n529), .ZN(new_n674));
  INV_X1    g0474(.A(new_n551), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n560), .A2(new_n561), .ZN(new_n676));
  OAI21_X1  g0476(.A(G169), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n567), .A2(G179), .A3(new_n551), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(new_n576), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n286), .A2(new_n327), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT94), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n304), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n301), .A2(KEYINPUT94), .A3(new_n303), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(G169), .B1(new_n688), .B2(new_n325), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n316), .A2(new_n321), .A3(new_n318), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n686), .B2(new_n687), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT95), .B1(new_n692), .B2(new_n503), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n309), .A2(new_n315), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n694), .A2(new_n320), .B1(new_n346), .B2(new_n317), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n301), .A2(KEYINPUT94), .A3(new_n303), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT94), .B1(new_n301), .B2(new_n303), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n316), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(G200), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n336), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n682), .A2(new_n683), .A3(new_n690), .A4(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n576), .B1(new_n677), .B2(new_n679), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n328), .A2(new_n338), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n705), .A3(new_n690), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n684), .A2(new_n689), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n699), .B1(new_n698), .B2(G200), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n294), .B(new_n332), .C1(new_n334), .C2(new_n322), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n707), .B1(new_n710), .B2(new_n700), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT96), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n602), .A2(new_n610), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n627), .A3(new_n657), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n503), .B1(new_n567), .B2(new_n551), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n544), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n677), .A2(new_n679), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n716), .A2(new_n578), .B1(new_n717), .B2(new_n544), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n660), .B2(new_n662), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n714), .A2(new_n718), .A3(new_n690), .A4(new_n701), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT96), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n706), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n673), .B1(new_n674), .B2(new_n724), .ZN(G369));
  NAND2_X1  g0525(.A1(new_n660), .A2(new_n662), .ZN(new_n726));
  INV_X1    g0526(.A(new_n256), .ZN(new_n727));
  OR3_X1    g0527(.A1(new_n727), .A2(KEYINPUT27), .A3(G20), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT27), .B1(new_n727), .B2(G20), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G213), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G343), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n732), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n714), .B1(new_n611), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n734), .A2(new_n639), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n720), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n656), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT98), .B(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n720), .A2(new_n734), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT99), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n735), .A2(new_n726), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n733), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n748), .ZN(G399));
  INV_X1    g0549(.A(new_n204), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G41), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n276), .A2(G116), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(G1), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n207), .B2(new_n752), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT101), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n722), .A2(KEYINPUT96), .ZN(new_n758));
  INV_X1    g0558(.A(new_n721), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n719), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n702), .A2(new_n690), .A3(new_n705), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n732), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n757), .B1(new_n762), .B2(KEYINPUT29), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  OAI211_X1 g0564(.A(KEYINPUT101), .B(new_n764), .C1(new_n724), .C2(new_n732), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n682), .A2(new_n690), .A3(new_n701), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT26), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n690), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n722), .A2(new_n721), .B1(KEYINPUT26), .B2(new_n704), .ZN(new_n769));
  OAI211_X1 g0569(.A(KEYINPUT29), .B(new_n734), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n628), .A2(new_n663), .A3(new_n339), .A4(new_n734), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n648), .A2(G179), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n773), .A2(new_n618), .A3(new_n698), .A4(new_n562), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n562), .A2(new_n322), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n616), .A2(new_n617), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n647), .A2(new_n777), .A3(new_n326), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n775), .B(KEYINPUT30), .C1(new_n776), .C2(new_n778), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n732), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT31), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(KEYINPUT31), .B(new_n732), .C1(new_n781), .C2(new_n782), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n772), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n740), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n771), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n756), .B1(new_n789), .B2(G1), .ZN(G364));
  NOR2_X1   g0590(.A1(new_n244), .A2(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n313), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n751), .A2(new_n793), .A3(KEYINPUT102), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT102), .B1(new_n751), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n742), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n740), .B2(new_n739), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n209), .B1(G20), .B2(new_n323), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n210), .A2(new_n326), .A3(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n492), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n334), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n493), .A2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n267), .B(new_n807), .C1(G326), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n210), .A2(G179), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(new_n334), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n811), .A2(new_n334), .A3(new_n503), .ZN(new_n814));
  INV_X1    g0614(.A(G329), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT105), .Z(new_n817));
  NOR2_X1   g0617(.A1(new_n808), .A2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT33), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(G317), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(G317), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n210), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n811), .A2(G190), .A3(G200), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n825), .A2(G294), .B1(new_n827), .B2(G303), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n810), .A2(new_n817), .A3(new_n822), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n814), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G159), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  INV_X1    g0632(.A(new_n818), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n833), .A2(new_n454), .B1(new_n826), .B2(new_n275), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n824), .A2(new_n278), .ZN(new_n836));
  INV_X1    g0636(.A(G58), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n803), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(G50), .C2(new_n809), .ZN(new_n839));
  INV_X1    g0639(.A(new_n812), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n471), .B1(new_n840), .B2(G107), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n806), .A2(KEYINPUT104), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n806), .A2(KEYINPUT104), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G77), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n835), .A2(new_n839), .A3(new_n841), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n801), .B1(new_n829), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(G13), .A2(G33), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(G20), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n800), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n482), .A2(new_n483), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n750), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n310), .B2(new_n208), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n237), .B2(new_n310), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n267), .A2(new_n204), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT103), .Z(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(G355), .B1(new_n300), .B2(new_n750), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n853), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n848), .A2(new_n862), .A3(new_n796), .ZN(new_n863));
  INV_X1    g0663(.A(new_n851), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n739), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n799), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G396));
  NAND2_X1  g0667(.A1(new_n760), .A2(new_n761), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n412), .A2(new_n732), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n420), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n416), .A2(new_n419), .A3(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT107), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n868), .A2(new_n734), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n668), .A2(new_n732), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n762), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n797), .B1(new_n878), .B2(new_n788), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n788), .B2(new_n878), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n801), .A2(new_n850), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n797), .B1(G77), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n833), .A2(KEYINPUT106), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n833), .A2(KEYINPUT106), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n845), .A2(G116), .B1(new_n886), .B2(G283), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n812), .A2(new_n275), .ZN(new_n888));
  INV_X1    g0688(.A(G294), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n803), .A2(new_n889), .B1(new_n389), .B2(new_n826), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n888), .B(new_n890), .C1(G303), .C2(new_n809), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n267), .B(new_n836), .C1(G311), .C2(new_n830), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n803), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(G143), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n809), .A2(G137), .B1(G150), .B2(new_n818), .ZN(new_n896));
  INV_X1    g0696(.A(G159), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n895), .B(new_n896), .C1(new_n844), .C2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT34), .Z(new_n899));
  INV_X1    g0699(.A(new_n854), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(G132), .B2(new_n830), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n825), .A2(G58), .B1(new_n840), .B2(G68), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n901), .B(new_n902), .C1(new_n373), .C2(new_n826), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n893), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n882), .B1(new_n904), .B2(new_n800), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n877), .B2(new_n850), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n880), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(G384));
  OR2_X1    g0708(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(G116), .A4(new_n211), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT36), .Z(new_n912));
  OAI211_X1 g0712(.A(new_n208), .B(G77), .C1(new_n837), .C2(new_n454), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n373), .A2(G68), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n313), .B(G13), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n460), .A2(new_n734), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n465), .B(new_n918), .C1(new_n448), .C2(new_n460), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n437), .A2(new_n440), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n446), .B1(new_n445), .B2(KEYINPUT14), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n442), .A2(KEYINPUT74), .A3(new_n443), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT108), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n917), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT108), .B1(new_n448), .B2(new_n918), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n787), .A3(new_n877), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT38), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n477), .B1(new_n485), .B2(new_n454), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n479), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n361), .A3(new_n486), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n469), .ZN(new_n934));
  INV_X1    g0734(.A(new_n730), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n521), .A2(new_n526), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n670), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n523), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n936), .A3(new_n510), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n487), .A2(new_n518), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n487), .B2(new_n506), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n487), .A2(new_n730), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT37), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n940), .A2(KEYINPUT37), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n930), .B1(new_n938), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(KEYINPUT37), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n944), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(KEYINPUT38), .C1(new_n527), .C2(new_n936), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT110), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n927), .A2(new_n787), .A3(new_n952), .A4(new_n877), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n929), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT40), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n522), .A2(new_n935), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n942), .A2(KEYINPUT109), .A3(KEYINPUT37), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n524), .A2(new_n957), .A3(new_n510), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT37), .B1(new_n943), .B2(KEYINPUT109), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n507), .A2(new_n508), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n957), .B1(new_n667), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n930), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n950), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n927), .A2(new_n787), .A3(KEYINPUT40), .A4(new_n877), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n956), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n529), .A2(new_n787), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n971), .A2(new_n740), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n763), .A2(new_n765), .A3(new_n529), .A4(new_n770), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n673), .ZN(new_n975));
  INV_X1    g0775(.A(new_n927), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n416), .A2(new_n732), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n875), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n951), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT39), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n966), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n462), .A2(new_n732), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n946), .A2(KEYINPUT39), .A3(new_n950), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n666), .A2(new_n519), .A3(new_n730), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n975), .B(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n973), .A2(new_n988), .B1(new_n313), .B2(new_n791), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n973), .A2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n916), .B1(new_n989), .B2(new_n990), .ZN(G367));
  NAND2_X1  g0791(.A1(new_n333), .A2(new_n732), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n711), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n690), .B2(new_n992), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(new_n864), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n852), .B1(new_n204), .B2(new_n247), .C1(new_n856), .C2(new_n228), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n797), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n824), .A2(new_n389), .ZN(new_n998));
  INV_X1    g0798(.A(G303), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n803), .A2(new_n999), .B1(new_n278), .B2(new_n812), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(G311), .C2(new_n809), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n813), .B2(new_n844), .C1(new_n889), .C2(new_n885), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n854), .B1(G317), .B2(new_n830), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n826), .B2(new_n300), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n267), .B1(new_n814), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n809), .B2(G143), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n894), .A2(G150), .B1(G68), .B2(new_n825), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n827), .A2(G58), .B1(new_n840), .B2(G77), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n844), .A2(new_n373), .B1(new_n885), .B2(new_n897), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1002), .A2(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n997), .B1(new_n1016), .B2(new_n800), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n995), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n682), .A2(new_n732), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n718), .B1(new_n576), .B2(new_n734), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n748), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT45), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n748), .A2(new_n1021), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT44), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n743), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1023), .A2(new_n743), .A3(new_n1025), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n736), .B(new_n746), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT113), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n741), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n741), .B(new_n1032), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n789), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n751), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n793), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT112), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1021), .B(KEYINPUT111), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1027), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT112), .B1(new_n1046), .B2(new_n743), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n736), .A2(new_n746), .A3(new_n1021), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT42), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n726), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n703), .B1(new_n1047), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1054), .B(new_n1055), .C1(new_n1057), .C2(new_n732), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1048), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1059));
  AND4_X1   g0859(.A1(new_n1042), .A2(new_n1051), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1051), .A2(new_n1059), .B1(new_n1058), .B2(new_n1042), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1018), .B1(new_n1041), .B2(new_n1062), .ZN(G387));
  OAI211_X1 g0863(.A(new_n753), .B(new_n310), .C1(new_n454), .C2(new_n342), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(KEYINPUT114), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n363), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n363), .B2(G50), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1068), .C1(new_n1064), .C2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n855), .B1(new_n1066), .B2(new_n1070), .C1(new_n225), .C2(new_n310), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n860), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(G107), .B2(new_n204), .C1(new_n753), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n852), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n797), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n736), .A2(new_n864), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n803), .A2(new_n373), .B1(new_n454), .B2(new_n806), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n363), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n818), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n900), .B1(G150), .B2(new_n830), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n825), .A2(new_n248), .B1(new_n840), .B2(G97), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n809), .A2(G159), .B1(G77), .B2(new_n827), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n854), .B1(G326), .B2(new_n830), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n824), .A2(new_n813), .B1(new_n826), .B2(new_n889), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G322), .A2(new_n809), .B1(new_n894), .B2(G317), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n805), .B2(new_n885), .C1(new_n999), .C2(new_n844), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1084), .B1(new_n300), .B2(new_n812), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1075), .B(new_n1076), .C1(new_n800), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1036), .B2(new_n793), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n789), .A2(new_n1036), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n751), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n789), .A2(new_n1036), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  INV_X1    g0900(.A(new_n1029), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n743), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n771), .A2(new_n788), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1037), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1030), .A2(new_n1097), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n751), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n793), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G68), .A2(new_n827), .B1(new_n830), .B2(G143), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n886), .A2(G50), .B1(KEYINPUT115), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(KEYINPUT115), .B2(new_n1110), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G150), .A2(new_n809), .B1(new_n894), .B2(G159), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n888), .B(new_n900), .C1(G77), .C2(new_n825), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n363), .B2(new_n844), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n806), .A2(new_n889), .B1(new_n826), .B2(new_n813), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n471), .B1(new_n814), .B2(new_n804), .C1(new_n389), .C2(new_n812), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(G116), .C2(new_n825), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n999), .B2(new_n885), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G317), .A2(new_n809), .B1(new_n894), .B2(G311), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT52), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n800), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n233), .A2(new_n856), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n853), .B1(G97), .B2(new_n750), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n796), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1125), .B(new_n1129), .C1(new_n1047), .C2(new_n864), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1108), .A2(new_n1109), .A3(new_n1130), .ZN(G390));
  OAI211_X1 g0931(.A(new_n734), .B(new_n874), .C1(new_n768), .C2(new_n769), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n978), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n927), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n983), .B1(new_n950), .B2(new_n965), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n927), .A2(new_n787), .A3(new_n740), .A4(new_n877), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n875), .A2(new_n978), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n983), .B1(new_n1138), .B2(new_n927), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT39), .B1(new_n950), .B2(new_n965), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n946), .A2(new_n950), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(KEYINPUT39), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1136), .B(new_n1137), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1135), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n976), .B1(new_n1132), .B2(new_n978), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n983), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n977), .B1(new_n762), .B2(new_n874), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n976), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n982), .A2(new_n984), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n927), .A2(new_n787), .A3(G330), .A4(new_n877), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(new_n792), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n849), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n809), .A2(G128), .ZN(new_n1156));
  OR3_X1    g0956(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n365), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT53), .B1(new_n826), .B2(new_n365), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n471), .B1(new_n830), .B2(G125), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n894), .A2(G132), .B1(G159), .B2(new_n825), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n373), .B2(new_n812), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n844), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n885), .A2(new_n1008), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1160), .A2(new_n1162), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n825), .A2(G77), .B1(new_n840), .B2(G68), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n809), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1167), .B1(new_n300), .B2(new_n803), .C1(new_n1168), .C2(new_n813), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n844), .A2(new_n278), .B1(new_n885), .B2(new_n389), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n471), .B1(new_n814), .B2(new_n889), .C1(new_n275), .C2(new_n826), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n800), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n797), .C1(new_n1078), .C2(new_n881), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT117), .Z(new_n1175));
  AOI21_X1  g0975(.A(new_n1154), .B1(new_n1155), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n787), .A2(new_n740), .A3(new_n877), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n976), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1152), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1138), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n787), .A2(G330), .A3(new_n877), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n976), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n978), .A3(new_n1132), .A4(new_n1137), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n529), .A2(G330), .A3(new_n787), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1184), .A2(new_n673), .A3(new_n974), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n752), .B1(new_n1153), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1152), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n872), .B(new_n869), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n732), .B(new_n1189), .C1(new_n760), .C2(new_n761), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n927), .B1(new_n1190), .B2(new_n977), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(new_n1147), .B1(new_n982), .B2(new_n984), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1188), .B1(new_n1192), .B2(new_n1146), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n974), .A2(new_n673), .A3(new_n1185), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1137), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n1133), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1196), .A2(new_n1182), .B1(new_n1179), .B2(new_n1138), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n1198), .A3(new_n1143), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT116), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  AOI221_X4 g1000(.A(new_n1195), .B1(new_n1134), .B2(new_n1135), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1150), .B1(new_n979), .B2(new_n983), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1152), .B1(new_n1202), .B2(new_n1136), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1186), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AND4_X1   g1004(.A1(KEYINPUT116), .A2(new_n1204), .A3(new_n1199), .A4(new_n751), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1176), .B1(new_n1200), .B2(new_n1205), .ZN(G378));
  INV_X1    g1006(.A(new_n987), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n928), .A2(KEYINPUT110), .B1(new_n946), .B2(new_n950), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT40), .B1(new_n1208), .B2(new_n953), .ZN(new_n1209));
  OAI21_X1  g1009(.A(G330), .B1(new_n967), .B2(new_n968), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n386), .A2(new_n423), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n378), .A2(new_n935), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1212), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n386), .A2(new_n423), .A3(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1216), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1214), .B1(new_n386), .B2(new_n423), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n665), .B(new_n1212), .C1(new_n382), .C2(new_n385), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1209), .A2(new_n1210), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1222), .ZN(new_n1224));
  INV_X1    g1024(.A(G330), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n968), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n966), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n956), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1207), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n956), .A2(new_n1227), .A3(new_n1224), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n987), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(KEYINPUT120), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1194), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1153), .B2(new_n1197), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT120), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n1207), .C1(new_n1223), .C2(new_n1228), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n752), .B1(new_n1241), .B2(new_n1235), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1233), .A2(new_n793), .A3(new_n1237), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n797), .B1(G50), .B2(new_n881), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n814), .A2(new_n813), .B1(new_n826), .B2(new_n342), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n900), .A2(new_n553), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(G58), .C2(new_n840), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT118), .Z(new_n1249));
  AOI22_X1  g1049(.A1(new_n809), .A2(G116), .B1(G68), .B2(new_n825), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT119), .Z(new_n1251));
  OAI22_X1  g1051(.A1(new_n803), .A2(new_n389), .B1(new_n278), .B2(new_n833), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n806), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n248), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT58), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n809), .A2(G125), .B1(new_n1253), .B2(G137), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1163), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n825), .A2(G150), .B1(new_n827), .B2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n894), .A2(G128), .B1(G132), .B2(new_n818), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G33), .A2(G41), .ZN(new_n1265));
  INV_X1    g1065(.A(G124), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1265), .B1(new_n814), .B2(new_n1266), .C1(new_n897), .C2(new_n812), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1263), .B2(KEYINPUT59), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1265), .A2(G50), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1264), .A2(new_n1268), .B1(new_n1247), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1257), .A2(new_n1258), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1245), .B1(new_n1271), .B2(new_n800), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1222), .B2(new_n850), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1244), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1243), .A2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n976), .A2(new_n849), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT121), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n809), .A2(G132), .B1(G159), .B2(new_n827), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n1278), .B1(new_n373), .B2(new_n824), .C1(new_n1008), .C2(new_n803), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n900), .B1(G128), .B2(new_n830), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n837), .B2(new_n812), .C1(new_n365), .C2(new_n806), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n886), .A2(new_n1260), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n845), .A2(G107), .B1(new_n886), .B2(G116), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n1168), .A2(new_n889), .B1(new_n278), .B2(new_n826), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n803), .A2(new_n813), .B1(new_n247), .B2(new_n824), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n471), .B1(new_n814), .B2(new_n999), .C1(new_n342), .C2(new_n812), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1282), .A2(new_n1283), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n797), .B1(G68), .B2(new_n881), .C1(new_n1289), .C2(new_n801), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1197), .A2(new_n792), .B1(new_n1277), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1198), .A2(new_n1039), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(G381));
  INV_X1    g1095(.A(G375), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1104), .B1(new_n1103), .B2(new_n1036), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n792), .B1(new_n1297), .B2(new_n1039), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1298), .A2(new_n1299), .B1(new_n995), .B2(new_n1017), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n866), .B(new_n1096), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1187), .A2(new_n1199), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1176), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1296), .A2(new_n1300), .A3(new_n1302), .A4(new_n1304), .ZN(G407));
  INV_X1    g1105(.A(G213), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G343), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1296), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  NAND2_X1  g1109(.A1(G393), .A2(G396), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1301), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(KEYINPUT123), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT124), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(G390), .A3(new_n1314), .A4(new_n1018), .ZN(new_n1315));
  INV_X1    g1115(.A(G390), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G387), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1300), .B2(G390), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT123), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1311), .B(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1316), .B2(G387), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1300), .A2(KEYINPUT125), .A3(G390), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1322), .A2(new_n1324), .A3(new_n1317), .A4(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1320), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1243), .A2(G378), .A3(new_n1274), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n793), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1273), .B(new_n1331), .C1(new_n1238), .C2(new_n1039), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1304), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1307), .B1(new_n1329), .B2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1194), .A2(new_n1197), .A3(KEYINPUT60), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1335), .A2(new_n751), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT60), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1293), .B1(new_n1198), .B2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1291), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(G384), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1339), .A2(G384), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1307), .ZN(new_n1343));
  INV_X1    g1143(.A(G2897), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OR3_X1    g1145(.A1(new_n1341), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1345), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1328), .B1(new_n1334), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(KEYINPUT126), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT126), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1351), .B(new_n1328), .C1(new_n1334), .C2(new_n1348), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1334), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(KEYINPUT62), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1350), .A2(new_n1352), .A3(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT122), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1354), .A2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1334), .A2(KEYINPUT122), .A3(new_n1353), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT62), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1327), .B1(new_n1356), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1358), .A2(new_n1362), .A3(new_n1359), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1320), .A2(new_n1326), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1349), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1363), .A2(new_n1364), .A3(new_n1365), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1361), .A2(new_n1367), .ZN(G405));
  OAI21_X1  g1168(.A(KEYINPUT127), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1327), .A2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(G375), .A2(new_n1304), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT127), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1353), .A2(new_n1372), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1371), .A2(new_n1329), .A3(new_n1373), .ZN(new_n1374));
  AND3_X1   g1174(.A1(new_n1320), .A2(new_n1326), .A3(new_n1369), .ZN(new_n1375));
  OR3_X1    g1175(.A1(new_n1370), .A2(new_n1374), .A3(new_n1375), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1374), .B1(new_n1370), .B2(new_n1375), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(G402));
endmodule


