//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n213), .B(new_n224), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n215), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n245), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G179), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n206), .A2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT5), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT76), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n260), .B2(KEYINPUT5), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n254), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT76), .B1(new_n256), .B2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n257), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(new_n262), .B2(KEYINPUT76), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  INV_X1    g0071(.A(new_n225), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n264), .A2(G257), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(G244), .A4(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT4), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G283), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n229), .A2(new_n253), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n288), .A2(KEYINPUT75), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT75), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n252), .B(new_n275), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT77), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n227), .A2(new_n228), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n284), .A2(new_n296), .A3(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n277), .A2(new_n279), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT7), .B1(new_n298), .B2(new_n207), .ZN(new_n299));
  OAI21_X1  g0099(.A(G107), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT6), .ZN(new_n301));
  INV_X1    g0101(.A(G97), .ZN(new_n302));
  INV_X1    g0102(.A(G107), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G97), .A2(G107), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n303), .A2(KEYINPUT73), .A3(KEYINPUT6), .A4(G97), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT6), .A2(G97), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(G107), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G77), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(KEYINPUT72), .A3(G77), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n311), .A2(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n300), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n311), .A2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n317), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n321), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n295), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G97), .ZN(new_n326));
  INV_X1    g0126(.A(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n295), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n206), .A2(G33), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(G97), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n288), .A2(new_n289), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n275), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n324), .A2(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n275), .B1(new_n290), .B2(new_n291), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n333), .A2(new_n275), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G190), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n324), .A2(new_n339), .A3(new_n331), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n293), .A2(new_n335), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(G1), .B1(new_n260), .B2(new_n267), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n274), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G226), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n254), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n284), .A2(G222), .A3(new_n280), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n284), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n346), .B1(new_n315), .B2(new_n284), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI211_X1 g0149(.A(new_n343), .B(new_n345), .C1(new_n349), .C2(new_n289), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n350), .A2(new_n252), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n206), .A2(G20), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n328), .A2(G50), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT8), .B(G58), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n207), .A2(G33), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n354), .A2(new_n355), .B1(new_n356), .B2(new_n314), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G20), .B2(new_n203), .ZN(new_n358));
  INV_X1    g0158(.A(new_n295), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n353), .B1(G50), .B2(new_n325), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n350), .B2(G169), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(G190), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n350), .A2(new_n367), .B1(new_n360), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n362), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT67), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n354), .A2(new_n314), .B1(new_n207), .B2(new_n315), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n355), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n295), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT66), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n315), .B1(new_n206), .B2(G20), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n328), .A2(new_n381), .B1(new_n315), .B2(new_n327), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n347), .A2(new_n216), .B1(new_n303), .B2(new_n284), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n298), .A2(new_n235), .A3(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n289), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n254), .A2(new_n342), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n343), .B1(G244), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(G169), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n375), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n252), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n380), .A2(new_n382), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(KEYINPUT67), .C1(G169), .C2(new_n389), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n389), .A2(G190), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n383), .B(new_n396), .C1(new_n367), .C2(new_n389), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n374), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n354), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n352), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n328), .B1(new_n327), .B2(new_n354), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT70), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT70), .B1(new_n277), .B2(new_n279), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n407), .B2(new_n207), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT71), .B(G68), .C1(new_n408), .C2(new_n297), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT70), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n278), .A2(G33), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT70), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n207), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n297), .B1(new_n416), .B2(new_n296), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n410), .B1(new_n417), .B2(new_n215), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G58), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(new_n215), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(new_n201), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(G20), .B1(G159), .B2(new_n313), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT16), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n359), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n297), .B2(new_n299), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n427), .B2(new_n423), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n404), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n284), .A2(new_n280), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n347), .B2(new_n344), .C1(new_n348), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n289), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n343), .B1(G232), .B2(new_n387), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n332), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(G179), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT18), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n297), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n405), .A2(new_n406), .A3(G20), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(KEYINPUT7), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT71), .B1(new_n442), .B2(G68), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n417), .A2(new_n410), .A3(new_n215), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n425), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n295), .A3(new_n429), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n434), .A2(new_n447), .A3(new_n435), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n437), .B2(G200), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n403), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n438), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n424), .B1(new_n409), .B2(new_n418), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n455), .A2(new_n359), .A3(new_n428), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n453), .B(new_n454), .C1(new_n456), .C2(new_n404), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n446), .A2(KEYINPUT17), .A3(new_n403), .A4(new_n449), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n439), .A2(new_n452), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n432), .B2(new_n344), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n298), .A2(new_n235), .A3(new_n280), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n289), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n343), .B1(G238), .B2(new_n387), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT13), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT13), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(G190), .A3(new_n468), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n314), .A2(new_n202), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n355), .A2(new_n315), .B1(new_n207), .B2(G68), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n295), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT11), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n325), .A2(G68), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT12), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT68), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n328), .A2(G68), .A3(new_n352), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n475), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n470), .A2(new_n471), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT69), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT69), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n470), .A2(new_n471), .A3(new_n488), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT14), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n469), .A2(new_n491), .A3(G169), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n252), .B2(new_n469), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n469), .B2(G169), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n484), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n399), .A2(new_n459), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n207), .B2(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n303), .A2(KEYINPUT23), .A3(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n277), .A2(new_n279), .A3(new_n207), .A4(G87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n284), .A2(new_n506), .A3(new_n207), .A4(G87), .ZN(new_n507));
  AOI211_X1 g0307(.A(KEYINPUT24), .B(new_n503), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n507), .ZN(new_n510));
  INV_X1    g0310(.A(new_n503), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n295), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n284), .A2(G257), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G294), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n277), .A2(new_n279), .A3(G250), .A4(new_n280), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n289), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n270), .A2(new_n274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n264), .A2(G264), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT25), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n325), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n327), .A2(KEYINPUT25), .A3(new_n303), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n330), .A2(G107), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n517), .A2(new_n289), .B1(new_n264), .B2(G264), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G190), .A3(new_n519), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n513), .A2(new_n522), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT86), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n521), .A2(new_n532), .A3(G169), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n531), .B(new_n533), .C1(new_n252), .C2(new_n521), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n513), .A2(new_n526), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT20), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(G33), .B2(G283), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n276), .A2(G97), .ZN(new_n540));
  INV_X1    g0340(.A(G116), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n539), .A2(new_n540), .B1(G20), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n542), .B2(new_n295), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n328), .A2(G116), .A3(new_n329), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n327), .A2(new_n541), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n542), .A2(new_n295), .A3(KEYINPUT82), .A4(new_n537), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n277), .A2(new_n279), .A3(G264), .A4(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n277), .A2(new_n279), .A3(G257), .A4(new_n280), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT81), .B(G303), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n284), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n289), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n264), .A2(G270), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n519), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n550), .B(KEYINPUT85), .C1(new_n558), .C2(new_n367), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n264), .A2(G270), .B1(new_n270), .B2(new_n274), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n367), .B1(new_n561), .B2(new_n555), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n562), .B2(new_n549), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(G190), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n549), .A2(new_n557), .A3(G169), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n549), .A2(new_n557), .A3(new_n568), .A4(G169), .ZN(new_n569));
  XOR2_X1   g0369(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n557), .A2(KEYINPUT21), .A3(G169), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n557), .A2(new_n252), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n549), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n565), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n254), .A2(new_n218), .A3(new_n268), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n274), .A2(KEYINPUT78), .A3(new_n268), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT78), .ZN(new_n578));
  OAI21_X1  g0378(.A(G274), .B1(new_n253), .B2(new_n225), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n255), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n277), .A2(new_n279), .A3(G244), .A4(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n277), .A2(new_n279), .A3(G238), .A4(new_n280), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n276), .C2(new_n541), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n289), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n585), .A3(G190), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n284), .A2(new_n207), .A3(G68), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n207), .B1(new_n460), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n305), .A2(new_n217), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n355), .B2(new_n302), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n295), .B1(new_n327), .B2(new_n377), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n330), .A2(G87), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n587), .A2(new_n588), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n581), .A2(new_n585), .A3(new_n252), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(KEYINPUT79), .ZN(new_n600));
  INV_X1    g0400(.A(new_n377), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n330), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT80), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(KEYINPUT79), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n596), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(KEYINPUT80), .B1(new_n332), .B2(new_n586), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n598), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n575), .A2(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n341), .A2(new_n497), .A3(new_n536), .A4(new_n611), .ZN(G372));
  AND3_X1   g0412(.A1(new_n439), .A2(KEYINPUT89), .A3(new_n457), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT89), .B1(new_n439), .B2(new_n457), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n495), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n395), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n391), .A2(KEYINPUT90), .A3(new_n392), .A4(new_n394), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n616), .B1(new_n621), .B2(new_n490), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n452), .A2(new_n458), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n373), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n369), .A2(new_n372), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n362), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n586), .A2(new_n332), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n607), .A3(new_n599), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n598), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n632), .B(new_n335), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n335), .B1(new_n633), .B2(new_n634), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n610), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n635), .A2(KEYINPUT88), .A3(new_n636), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n340), .A2(new_n337), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n598), .A2(new_n631), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n529), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n640), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT87), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n640), .A2(new_n645), .A3(new_n650), .A4(new_n647), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n534), .A2(new_n535), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n571), .A2(new_n574), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n649), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n644), .A2(new_n655), .A3(new_n631), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n497), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n629), .A2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT91), .Z(new_n663));
  XNOR2_X1  g0463(.A(KEYINPUT92), .B(G343), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n652), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n665), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT94), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT94), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n652), .A2(new_n670), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n535), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT93), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n669), .A2(new_n671), .B1(new_n673), .B2(new_n536), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n653), .A2(new_n665), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n666), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n665), .A2(new_n550), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n653), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n575), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n676), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n210), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n592), .A2(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n231), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n656), .A2(new_n690), .A3(new_n665), .ZN(new_n691));
  MUX2_X1   g0491(.A(new_n635), .B(new_n641), .S(new_n636), .Z(new_n692));
  NOR2_X1   g0492(.A1(new_n652), .A2(new_n653), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n631), .B1(new_n693), .B2(new_n648), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n665), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n581), .A2(new_n585), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n275), .A3(new_n333), .A4(new_n527), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n558), .A2(G179), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n699), .A2(G179), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n336), .A2(new_n703), .A3(new_n521), .A4(new_n557), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n518), .A2(new_n520), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n586), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n573), .A3(new_n338), .A4(KEYINPUT30), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT31), .B1(new_n708), .B2(new_n667), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n334), .A2(new_n705), .A3(new_n586), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT30), .B1(new_n711), .B2(new_n573), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n521), .A2(new_n557), .A3(new_n586), .A4(new_n252), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT75), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n333), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n288), .A2(KEYINPUT75), .A3(new_n289), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n275), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n710), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT95), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n707), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n667), .A2(KEYINPUT31), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n709), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n611), .A2(new_n341), .A3(new_n536), .A4(new_n665), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n728), .A3(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n697), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n689), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n680), .ZN(new_n733));
  INV_X1    g0533(.A(G13), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n206), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n684), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n679), .ZN(new_n740));
  INV_X1    g0540(.A(new_n738), .ZN(new_n741));
  INV_X1    g0541(.A(new_n229), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n207), .B2(G169), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT97), .ZN(new_n744));
  NAND2_X1  g0544(.A1(G20), .A2(G179), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(G317), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT33), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n749), .A2(KEYINPUT33), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n447), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n207), .ZN(new_n755));
  INV_X1    g0555(.A(G303), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n207), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n752), .B1(new_n753), .B2(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n284), .B1(new_n762), .B2(G329), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(new_n760), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n745), .A2(new_n447), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n763), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n747), .A2(new_n447), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n207), .A2(new_n367), .A3(G179), .A4(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n759), .A2(new_n769), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n758), .A2(new_n217), .ZN(new_n778));
  INV_X1    g0578(.A(new_n748), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n215), .B1(new_n774), .B2(new_n303), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G50), .C2(new_n770), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n762), .A2(G159), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT32), .ZN(new_n783));
  INV_X1    g0583(.A(new_n755), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n782), .A2(KEYINPUT32), .B1(new_n784), .B2(G97), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n284), .B1(new_n768), .B2(new_n420), .ZN(new_n786));
  INV_X1    g0586(.A(new_n765), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G77), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n781), .A2(new_n783), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n744), .B1(new_n777), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n744), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT98), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n210), .A2(G355), .A3(new_n284), .ZN(new_n798));
  INV_X1    g0598(.A(new_n407), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n683), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n231), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n250), .A2(new_n267), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n798), .B1(G116), .B2(new_n210), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n741), .B(new_n790), .C1(new_n797), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n794), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n679), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n740), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  AND2_X1   g0608(.A1(new_n398), .A2(new_n665), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n656), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n667), .A2(new_n393), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n398), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n620), .B2(new_n812), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n656), .B2(new_n665), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n729), .B(new_n727), .C1(new_n811), .C2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n811), .A2(new_n815), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n738), .B1(new_n819), .B2(new_n730), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n787), .A2(G159), .B1(G143), .B2(new_n767), .ZN(new_n822));
  INV_X1    g0622(.A(new_n770), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n356), .C2(new_n779), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n407), .B1(G132), .B2(new_n762), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n758), .A2(new_n202), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n774), .A2(new_n215), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G58), .C2(new_n784), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n772), .A2(new_n779), .B1(new_n823), .B2(new_n756), .ZN(new_n834));
  INV_X1    g0634(.A(new_n758), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(G107), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n784), .A2(G97), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n768), .A2(new_n753), .B1(new_n761), .B2(new_n764), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n284), .B(new_n838), .C1(G116), .C2(new_n787), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n773), .A2(G87), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n836), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n744), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n744), .A2(new_n793), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT100), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n741), .B(new_n842), .C1(new_n845), .C2(new_n315), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n814), .B2(new_n793), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n821), .A2(new_n847), .ZN(G384));
  NOR2_X1   g0648(.A1(new_n735), .A2(new_n206), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT103), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n423), .B1(new_n443), .B2(new_n444), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT16), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n404), .B1(new_n853), .B2(new_n426), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n450), .B1(new_n854), .B2(new_n438), .ZN(new_n855));
  INV_X1    g0655(.A(new_n663), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n446), .A2(new_n403), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n453), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n663), .B1(new_n456), .B2(new_n404), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n450), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n858), .A2(new_n863), .B1(new_n459), .B2(new_n857), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n850), .B1(new_n864), .B2(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n858), .A2(new_n863), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n459), .A2(new_n857), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n850), .A3(new_n869), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n864), .A2(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n860), .A2(new_n450), .A3(new_n862), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(new_n861), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n452), .B(new_n458), .C1(new_n613), .C2(new_n614), .ZN(new_n878));
  INV_X1    g0678(.A(new_n862), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n874), .B(new_n875), .C1(new_n880), .C2(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n616), .A2(new_n665), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n485), .A2(new_n665), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n496), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n886), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n490), .B2(new_n495), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n395), .A2(new_n667), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n810), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n872), .A3(new_n871), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n615), .A2(new_n663), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n697), .A2(new_n497), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n629), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(G330), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n814), .B1(new_n887), .B2(new_n889), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n709), .B1(new_n708), .B2(new_n722), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n724), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n871), .A2(new_n872), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n875), .B1(new_n880), .B2(KEYINPUT38), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n905), .A2(new_n911), .A3(new_n908), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n910), .A2(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n497), .A2(new_n907), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n904), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n849), .B1(new_n903), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n903), .B2(new_n917), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n311), .A2(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n311), .A2(KEYINPUT35), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(G116), .A3(new_n230), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  OAI21_X1  g0723(.A(G77), .B1(new_n420), .B2(new_n215), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n246), .B1(new_n924), .B2(new_n231), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n734), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n923), .A3(new_n926), .ZN(G367));
  NAND2_X1  g0727(.A1(new_n669), .A2(new_n671), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n673), .A2(new_n536), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n675), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n324), .A2(new_n331), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n341), .B1(new_n931), .B2(new_n665), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n293), .A2(new_n335), .A3(new_n667), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n652), .A2(new_n645), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n667), .B1(new_n937), .B2(new_n640), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n935), .B2(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n597), .A2(new_n596), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n667), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(new_n631), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n632), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n940), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n936), .A2(new_n939), .A3(new_n947), .A4(new_n946), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n681), .ZN(new_n953));
  INV_X1    g0753(.A(new_n934), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n952), .B(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n684), .B(KEYINPUT41), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n676), .A2(new_n954), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n676), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n930), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n963), .A2(KEYINPUT45), .A3(new_n666), .A4(new_n934), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n676), .B2(new_n954), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n681), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n674), .A2(new_n675), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(KEYINPUT104), .A3(new_n680), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n680), .B1(new_n970), .B2(KEYINPUT104), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n963), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n971), .A3(new_n930), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n962), .A2(new_n967), .A3(new_n953), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n969), .A2(new_n731), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n957), .B1(new_n979), .B2(new_n731), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n956), .B1(new_n980), .B2(new_n737), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n768), .A2(new_n356), .B1(new_n765), .B2(new_n202), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n298), .B(new_n982), .C1(G137), .C2(new_n762), .ZN(new_n983));
  INV_X1    g0783(.A(G159), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n779), .A2(new_n984), .B1(new_n758), .B2(new_n420), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n755), .A2(new_n215), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n770), .A2(G143), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n773), .A2(G77), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n983), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n823), .A2(new_n764), .B1(new_n303), .B2(new_n755), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G294), .B2(new_n748), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n762), .A2(G317), .ZN(new_n993));
  INV_X1    g0793(.A(new_n553), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n787), .A2(G283), .B1(new_n994), .B2(new_n767), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n799), .B1(G97), .B2(new_n773), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n993), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n758), .A2(new_n541), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT105), .Z(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT47), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT47), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n791), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n800), .A2(new_n241), .B1(new_n683), .B2(new_n601), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n741), .B1(new_n795), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(new_n805), .C2(new_n945), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n981), .A2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n977), .A2(new_n737), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n686), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n210), .A3(new_n284), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(G107), .B2(new_n210), .ZN(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n1010), .C1(G68), .C2(G77), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n354), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n683), .B(new_n799), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n238), .A2(G45), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n738), .B1(new_n796), .B2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n768), .A2(new_n202), .B1(new_n765), .B2(new_n215), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n762), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n407), .B1(G97), .B2(new_n773), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n784), .A2(new_n601), .B1(new_n770), .B2(G159), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n400), .A2(new_n748), .B1(new_n835), .B2(G77), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n799), .B1(G326), .B2(new_n762), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n755), .A2(new_n772), .B1(new_n758), .B2(new_n753), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n787), .A2(new_n994), .B1(G317), .B2(new_n767), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n823), .B2(new_n766), .C1(new_n764), .C2(new_n779), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1026), .B1(new_n541), .B2(new_n774), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1019), .B1(new_n1036), .B2(new_n791), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n674), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n805), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT106), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n977), .A2(new_n731), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n684), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n977), .A2(new_n731), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1009), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(G393));
  NAND3_X1  g0844(.A1(new_n969), .A2(new_n737), .A3(new_n978), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n800), .A2(new_n245), .B1(G97), .B2(new_n683), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n741), .B1(new_n795), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n298), .B1(new_n766), .B2(new_n761), .C1(new_n774), .C2(new_n303), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G283), .B2(new_n835), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT107), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n755), .A2(new_n541), .B1(new_n765), .B2(new_n753), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n767), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n994), .C2(new_n748), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G143), .A2(new_n762), .B1(new_n787), .B2(new_n400), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n799), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n779), .A2(new_n202), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n840), .B1(new_n215), .B2(new_n758), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n755), .A2(new_n315), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n770), .A2(G150), .B1(G159), .B2(new_n767), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  AOI22_X1  g0862(.A1(new_n1050), .A2(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1047), .B1(new_n744), .B2(new_n1063), .C1(new_n934), .C2(new_n805), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n969), .A2(new_n978), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(new_n1041), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n979), .A2(new_n684), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1045), .B(new_n1064), .C1(new_n1066), .C2(new_n1067), .ZN(G390));
  AOI21_X1  g0868(.A(new_n1059), .B1(G116), .B2(new_n767), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT110), .Z(new_n1070));
  OAI22_X1  g0870(.A1(new_n303), .A2(new_n779), .B1(new_n823), .B2(new_n772), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n298), .B1(new_n765), .B2(new_n302), .C1(new_n753), .C2(new_n761), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1071), .A2(new_n778), .A3(new_n831), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT54), .B(G143), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n748), .A2(G137), .B1(new_n787), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT109), .Z(new_n1078));
  INV_X1    g0878(.A(G125), .ZN(new_n1079));
  INV_X1    g0879(.A(G132), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n284), .B1(new_n761), .B2(new_n1079), .C1(new_n768), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT53), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n835), .B2(G150), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n356), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(G128), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n823), .A2(new_n1086), .B1(new_n774), .B2(new_n202), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G159), .B2(new_n784), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1078), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n744), .B1(new_n1074), .B2(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n741), .B(new_n1090), .C1(new_n845), .C2(new_n354), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n882), .B2(new_n793), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n893), .B1(new_n656), .B2(new_n809), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n883), .B1(new_n1093), .B2(new_n890), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n873), .A2(new_n881), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n814), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n891), .B1(new_n695), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n890), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n912), .A2(new_n1099), .A3(new_n883), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n905), .A2(new_n904), .A3(new_n908), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n730), .A2(new_n814), .A3(new_n1098), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1095), .A2(new_n1104), .A3(new_n1100), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1092), .B1(new_n1106), .B2(new_n736), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n908), .A2(new_n904), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n497), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n901), .A2(new_n629), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1093), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1098), .B1(new_n730), .B2(new_n814), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n1102), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1108), .A2(new_n814), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1114), .B2(new_n890), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1104), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1110), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1103), .A2(new_n1117), .A3(new_n1105), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n684), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1110), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT108), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT108), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1125), .A3(new_n1106), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1107), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n910), .A2(new_n911), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n360), .A2(new_n663), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n374), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n374), .A2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n374), .A2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n374), .A2(new_n1133), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1131), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1130), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1130), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n900), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1130), .A2(new_n1142), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n883), .B1(new_n873), .B2(new_n881), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n896), .A2(new_n898), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1130), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1129), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n685), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1145), .A2(new_n1153), .A3(KEYINPUT118), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT118), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1148), .A2(new_n1151), .A3(new_n1158), .A4(new_n1152), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1157), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1156), .B1(new_n1160), .B2(KEYINPUT57), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1141), .A2(new_n793), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(G33), .A2(G41), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G50), .B(new_n1163), .C1(new_n407), .C2(new_n260), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT111), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n774), .A2(new_n420), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n758), .A2(new_n315), .B1(new_n761), .B2(new_n772), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n799), .A2(new_n1166), .A3(G41), .A4(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT112), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n768), .A2(new_n303), .B1(new_n377), .B2(new_n765), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n302), .A2(new_n779), .B1(new_n823), .B2(new_n541), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1169), .A2(new_n986), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1165), .B1(new_n1172), .B2(KEYINPUT58), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT113), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n787), .A2(G137), .B1(G128), .B2(new_n767), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n758), .B2(new_n1075), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1079), .A2(new_n823), .B1(new_n779), .B2(new_n1080), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G150), .C2(new_n784), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT59), .Z(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT114), .ZN(new_n1180));
  OR2_X1    g0980(.A1(KEYINPUT115), .A2(G124), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(KEYINPUT115), .A2(G124), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n762), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n1163), .C1(new_n984), .C2(new_n774), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1179), .B2(KEYINPUT114), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1180), .A2(new_n1185), .B1(KEYINPUT58), .B2(new_n1172), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n744), .B1(new_n1174), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT116), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n738), .B1(new_n844), .B2(G50), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1162), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n737), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1161), .A2(new_n1192), .ZN(G375));
  NOR2_X1   g0993(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n957), .B(KEYINPUT119), .Z(new_n1196));
  NAND4_X1  g0996(.A1(new_n1123), .A2(new_n1195), .A3(new_n1125), .A4(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1098), .A2(new_n793), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n541), .A2(new_n779), .B1(new_n823), .B2(new_n753), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G97), .B2(new_n835), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n784), .A2(new_n601), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n768), .A2(new_n772), .B1(new_n765), .B2(new_n303), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n284), .B(new_n1202), .C1(G303), .C2(new_n762), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n989), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n755), .A2(new_n202), .B1(new_n765), .B2(new_n356), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT121), .Z(new_n1206));
  NOR2_X1   g1006(.A1(new_n758), .A2(new_n984), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1207), .B(new_n1166), .C1(new_n748), .C2(new_n1076), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n770), .A2(G132), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT120), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n768), .A2(new_n824), .B1(new_n761), .B2(new_n1086), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n407), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n744), .B1(new_n1204), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n741), .B(new_n1214), .C1(new_n845), .C2(new_n215), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT122), .Z(new_n1216));
  NOR2_X1   g1016(.A1(new_n1198), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1120), .B2(new_n737), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1197), .A2(new_n1218), .ZN(G381));
  NOR4_X1   g1019(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n981), .A3(new_n1007), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G378), .A2(G375), .A3(new_n1221), .A4(G381), .ZN(G407));
  INV_X1    g1022(.A(G213), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n664), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1127), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G375), .C2(new_n1225), .ZN(G409));
  XNOR2_X1  g1026(.A(G393), .B(new_n807), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G390), .A2(new_n981), .A3(new_n1007), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G390), .B1(new_n981), .B2(new_n1007), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1161), .A2(G378), .A3(new_n1192), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1157), .A2(new_n1155), .A3(new_n1159), .A4(new_n1196), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1190), .B1(new_n1239), .B2(new_n737), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1127), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1244), .A3(new_n1127), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1237), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1224), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1194), .A2(KEYINPUT60), .A3(new_n1122), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n684), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1194), .B1(KEYINPUT60), .B2(new_n1122), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1218), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1248), .B(G384), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G384), .A2(new_n1248), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(new_n1253), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G384), .A2(new_n1248), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n1251), .C2(new_n1250), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1246), .A2(new_n1247), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1247), .A4(new_n1259), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT62), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1259), .A2(G2897), .A3(new_n1224), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1224), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1254), .A2(new_n1258), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1236), .B1(new_n1264), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1236), .B2(KEYINPUT61), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1232), .A2(new_n1235), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1262), .A2(new_n1280), .A3(new_n1263), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1260), .A2(new_n1280), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1273), .A2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(G375), .A2(new_n1127), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1237), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(KEYINPUT127), .A3(new_n1237), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1259), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1286), .A2(new_n1287), .A3(new_n1254), .A4(new_n1258), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1236), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1292), .B(new_n1293), .ZN(G402));
endmodule


