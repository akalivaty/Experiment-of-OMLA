//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G43gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT83), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n210), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(new_n209), .B2(new_n211), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(new_n213), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NOR4_X1   g025(.A1(KEYINPUT86), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(new_n214), .B2(new_n215), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n207), .B1(new_n230), .B2(new_n212), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n204), .A2(KEYINPUT85), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G50gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n202), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n205), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n220), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n231), .A2(KEYINPUT87), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT87), .B1(new_n231), .B2(new_n238), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT17), .B(new_n226), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G15gat), .B(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT16), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(G1gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G1gat), .B2(new_n242), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n245), .B(G8gat), .Z(new_n246));
  OR2_X1    g045(.A1(new_n224), .A2(new_n213), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n220), .B1(new_n224), .B2(new_n213), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n206), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n223), .B(new_n228), .ZN(new_n251));
  INV_X1    g050(.A(new_n212), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n206), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n205), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT85), .B(G50gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n202), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n221), .B1(new_n256), .B2(KEYINPUT15), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n250), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT87), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n261));
  OAI211_X1 g060(.A(new_n241), .B(new_n246), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G229gat), .A2(G233gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n246), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n226), .B1(new_n239), .B2(new_n240), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT90), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT18), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT11), .B(G169gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G197gat), .ZN(new_n272));
  XOR2_X1   g071(.A(G113gat), .B(G141gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n262), .A2(KEYINPUT18), .A3(new_n263), .A4(new_n266), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT89), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n246), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n266), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n263), .B(KEYINPUT13), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n269), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT90), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n276), .A2(new_n278), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n262), .A2(new_n266), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n286), .A2(KEYINPUT89), .A3(KEYINPUT18), .A4(new_n263), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n283), .A3(new_n282), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n275), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G230gat), .ZN(new_n294));
  INV_X1    g093(.A(G233gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G99gat), .A2(G106gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT8), .ZN(new_n298));
  NAND2_X1  g097(.A1(G85gat), .A2(G92gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G85gat), .ZN(new_n302));
  INV_X1    g101(.A(G92gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n298), .A2(new_n301), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G99gat), .ZN(new_n308));
  INV_X1    g107(.A(G106gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(KEYINPUT96), .A3(new_n297), .ZN(new_n315));
  AOI22_X1  g114(.A1(KEYINPUT8), .A2(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n316));
  AND3_X1   g115(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n310), .A2(KEYINPUT96), .A3(new_n297), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT96), .B1(new_n310), .B2(new_n297), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n306), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G71gat), .A2(G78gat), .ZN(new_n326));
  OR2_X1    g125(.A1(G71gat), .A2(G78gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G57gat), .B(G64gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n328), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n329), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n325), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT98), .B1(new_n322), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n306), .B1(new_n323), .B2(new_n324), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n337), .A2(KEYINPUT97), .B1(new_n311), .B2(new_n307), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n330), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n338), .A2(new_n340), .A3(new_n341), .A4(new_n325), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344));
  INV_X1    g143(.A(new_n311), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n306), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n312), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n306), .A2(new_n345), .A3(KEYINPUT93), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n339), .A3(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n336), .A2(new_n342), .A3(new_n343), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT10), .A3(new_n340), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n296), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n342), .A3(new_n349), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n296), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G176gat), .B(G204gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT99), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(G120gat), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n355), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n293), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT21), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n246), .B1(new_n365), .B2(new_n339), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G183gat), .ZN(new_n367));
  INV_X1    g166(.A(G231gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n295), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n366), .B(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n295), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G127gat), .B(G155gat), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n377), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n339), .A2(new_n365), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n381), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n261), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n265), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n351), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n241), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT94), .ZN(new_n391));
  NAND2_X1  g190(.A1(G232gat), .A2(G233gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT91), .Z(new_n393));
  INV_X1    g192(.A(KEYINPUT41), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n265), .B2(new_n351), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n388), .A2(new_n397), .A3(new_n241), .A4(new_n389), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n391), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G190gat), .B(G218gat), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n391), .A2(new_n400), .A3(new_n396), .A4(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G134gat), .B(G162gat), .Z(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT92), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n393), .A2(new_n394), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n402), .A2(new_n411), .A3(new_n403), .A4(new_n408), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n386), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(G113gat), .B(G120gat), .Z(new_n416));
  XNOR2_X1  g215(.A(G127gat), .B(G134gat), .ZN(new_n417));
  OR2_X1    g216(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n418));
  NAND2_X1  g217(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT70), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G127gat), .B(G134gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(KEYINPUT1), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT76), .ZN(new_n429));
  INV_X1    g228(.A(G155gat), .ZN(new_n430));
  INV_X1    g229(.A(G162gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G141gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G148gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n359), .A2(G141gat), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n428), .A2(KEYINPUT2), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n429), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n428), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT77), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n434), .A2(new_n435), .B1(KEYINPUT2), .B2(new_n428), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n442), .A3(new_n428), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n422), .A2(new_n427), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n422), .A2(new_n427), .A3(new_n446), .A4(KEYINPUT4), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n445), .A2(KEYINPUT3), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n445), .A2(KEYINPUT3), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT78), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n422), .A2(new_n427), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n422), .B2(new_n427), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n453), .B(new_n455), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n452), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n427), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n422), .A2(new_n427), .A3(new_n456), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n446), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n447), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT5), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT0), .B(G57gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(G85gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n460), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n449), .A2(new_n450), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n453), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT5), .B1(new_n481), .B2(new_n452), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n473), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n474), .A4(new_n476), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G204gat), .ZN(new_n488));
  INV_X1    g287(.A(G197gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT22), .ZN(new_n491));
  INV_X1    g290(.A(G218gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n376), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G211gat), .B(G218gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n495), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G226gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n295), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT29), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT27), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G183gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT65), .B(G183gat), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT27), .ZN(new_n510));
  NOR2_X1   g309(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G169gat), .A2(G176gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT26), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT67), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G183gat), .A2(G190gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT28), .B1(new_n524), .B2(G190gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n512), .A2(new_n521), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT64), .B(G176gat), .ZN(new_n527));
  INV_X1    g326(.A(G169gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT23), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n522), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n534), .B(new_n535), .C1(G183gat), .C2(G190gat), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n531), .A2(new_n513), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n513), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(KEYINPUT23), .B2(new_n514), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT65), .B(G183gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(G190gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n535), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n532), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT25), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n526), .A2(new_n537), .A3(KEYINPUT75), .A4(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n504), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n545), .A2(new_n501), .A3(new_n295), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n500), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n502), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n545), .A2(new_n503), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n499), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G8gat), .B(G36gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G64gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n303), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n551), .A2(new_n558), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT30), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n563), .A3(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n487), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G22gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT29), .ZN(new_n569));
  INV_X1    g368(.A(new_n498), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n495), .B1(new_n490), .B2(new_n493), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT3), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n446), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n499), .B1(new_n569), .B2(new_n455), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n500), .B1(KEYINPUT29), .B2(new_n454), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT29), .B1(new_n497), .B2(new_n498), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n445), .B1(new_n578), .B2(KEYINPUT3), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n579), .A3(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G228gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n574), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G50gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n204), .B(new_n582), .C1(new_n574), .C2(new_n583), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G78gat), .B(G106gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(new_n587), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n566), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598));
  NAND2_X1  g397(.A1(G227gat), .A2(G233gat), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n537), .A2(new_n544), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(new_n422), .A3(new_n427), .A4(new_n526), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n545), .A2(new_n462), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n603), .B2(KEYINPUT33), .ZN(new_n604));
  INV_X1    g403(.A(new_n599), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n545), .A2(new_n462), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n545), .A2(new_n462), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(KEYINPUT71), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(KEYINPUT32), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT72), .B(G15gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n202), .ZN(new_n613));
  XOR2_X1   g412(.A(G71gat), .B(G99gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n604), .A2(new_n610), .A3(new_n611), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(KEYINPUT32), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n599), .A3(new_n602), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT73), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT34), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n619), .B2(new_n620), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n616), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(new_n616), .B2(new_n618), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n597), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n616), .A2(new_n618), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n616), .A2(new_n624), .A3(new_n618), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT36), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n551), .A2(KEYINPUT37), .A3(new_n554), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT81), .B1(new_n555), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT81), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n639), .B(new_n636), .C1(new_n551), .C2(new_n554), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n635), .B(new_n558), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT38), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n560), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n644), .B(new_n558), .C1(new_n638), .C2(new_n640), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n549), .A2(new_n500), .A3(new_n550), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n499), .B1(new_n552), .B2(new_n553), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n485), .B(new_n486), .C1(new_n645), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n595), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n452), .B1(new_n451), .B2(new_n459), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n473), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n465), .A2(new_n461), .A3(new_n466), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n656), .B2(new_n658), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n661), .A2(new_n564), .A3(new_n477), .A4(new_n562), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n652), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n596), .B(new_n634), .C1(new_n651), .C2(new_n663), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n485), .A2(new_n486), .B1(new_n564), .B2(new_n562), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n630), .A2(KEYINPUT82), .A3(new_n631), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT82), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n625), .B2(new_n626), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n665), .A2(new_n652), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT35), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n591), .B(new_n594), .C1(new_n625), .C2(new_n626), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n670), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n669), .A2(new_n670), .B1(new_n665), .B2(new_n672), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n364), .B(new_n415), .C1(new_n664), .C2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n487), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  INV_X1    g476(.A(new_n565), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT101), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(KEYINPUT42), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n679), .B(KEYINPUT100), .Z(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(G8gat), .ZN(new_n685));
  OAI221_X1 g484(.A(new_n682), .B1(KEYINPUT42), .B2(new_n681), .C1(new_n683), .C2(new_n685), .ZN(G1325gat));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n666), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(G15gat), .B1(new_n674), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n633), .A2(G15gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n674), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n595), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n664), .A2(new_n673), .ZN(new_n695));
  INV_X1    g494(.A(new_n414), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n414), .B1(new_n664), .B2(new_n673), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n386), .A2(new_n364), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n487), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n700), .A2(new_n703), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n218), .A3(new_n675), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n219), .A3(new_n678), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n705), .B2(new_n565), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  AND2_X1   g513(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n202), .A3(new_n688), .A4(new_n703), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT103), .Z(new_n717));
  NAND4_X1  g516(.A1(new_n699), .A2(new_n633), .A3(new_n701), .A4(new_n704), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n702), .A2(new_n595), .A3(new_n704), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n255), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n652), .A2(new_n255), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n728), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n724), .A2(new_n726), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n729), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n725), .B2(new_n255), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n724), .B1(new_n732), .B2(new_n727), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n733), .ZN(G1331gat));
  AOI21_X1  g533(.A(new_n415), .B1(new_n664), .B2(new_n673), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n293), .A2(new_n363), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n675), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n565), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  OR3_X1    g544(.A1(new_n737), .A2(G71gat), .A3(new_n687), .ZN(new_n746));
  OAI21_X1  g545(.A(G71gat), .B1(new_n737), .B2(new_n634), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g548(.A1(new_n737), .A2(new_n652), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(G78gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  NAND4_X1  g551(.A1(new_n699), .A2(new_n385), .A3(new_n701), .A4(new_n736), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(G85gat), .A3(new_n675), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n386), .A2(new_n293), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT51), .B1(new_n697), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n700), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(new_n675), .A3(new_n362), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n302), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT107), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n754), .A2(G92gat), .A3(new_n678), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n758), .A2(new_n362), .A3(new_n678), .A4(new_n760), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n303), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n753), .B2(new_n634), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n758), .A2(new_n760), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n308), .A3(new_n362), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n773), .B2(new_n687), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n776), .B(new_n771), .C1(new_n773), .C2(new_n687), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1338gat));
  OAI21_X1  g577(.A(G106gat), .B1(new_n753), .B2(new_n652), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n772), .A2(new_n309), .A3(new_n362), .A4(new_n595), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT109), .B(G106gat), .C1(new_n753), .C2(new_n652), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1339gat));
  AOI21_X1  g587(.A(new_n263), .B1(new_n262), .B2(new_n266), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n266), .A2(new_n279), .A3(new_n281), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n274), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n285), .A2(new_n793), .A3(new_n362), .ZN(new_n794));
  AND4_X1   g593(.A1(new_n282), .A2(new_n284), .A3(new_n287), .A4(new_n289), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n350), .A2(new_n352), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  INV_X1    g598(.A(new_n296), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n350), .A2(new_n296), .A3(new_n352), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n360), .B(new_n801), .C1(new_n803), .C2(new_n353), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n797), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n803), .A2(new_n353), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n361), .B1(new_n353), .B2(new_n799), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n804), .A2(new_n805), .B1(new_n355), .B2(new_n361), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n414), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n285), .A2(new_n793), .A3(new_n810), .A4(new_n811), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n414), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n385), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n386), .A2(new_n796), .A3(new_n363), .A4(new_n414), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n487), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n821), .A2(new_n565), .A3(new_n652), .A4(new_n688), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n796), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n487), .B(new_n671), .C1(new_n819), .C2(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n565), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(G113gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n826), .B2(new_n796), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n822), .B2(new_n363), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n825), .A2(G120gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n363), .ZN(G1341gat));
  INV_X1    g629(.A(new_n825), .ZN(new_n831));
  AOI21_X1  g630(.A(G127gat), .B1(new_n831), .B2(new_n386), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n822), .A2(new_n385), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(G127gat), .B2(new_n833), .ZN(G1342gat));
  NOR3_X1   g633(.A1(new_n825), .A2(G134gat), .A3(new_n414), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n822), .B2(new_n414), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G1343gat));
  NOR3_X1   g639(.A1(new_n633), .A2(new_n487), .A3(new_n678), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n816), .B1(new_n414), .B2(new_n813), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n386), .ZN(new_n845));
  INV_X1    g644(.A(new_n812), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n293), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n696), .B1(new_n847), .B2(new_n794), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT113), .B(new_n385), .C1(new_n848), .C2(new_n816), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n820), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n595), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n842), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n820), .B1(new_n844), .B2(new_n386), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n595), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(G141gat), .A3(new_n293), .A4(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n634), .A2(KEYINPUT114), .A3(new_n595), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n633), .B2(new_n652), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n821), .A2(new_n565), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n433), .B1(new_n862), .B2(new_n796), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(new_n862), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n359), .A3(new_n362), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n362), .A3(new_n855), .A4(new_n841), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n359), .A2(KEYINPUT59), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT116), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n385), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n820), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n652), .A2(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n853), .A2(new_n595), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT57), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n362), .A3(new_n841), .A4(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n359), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n880), .A2(new_n881), .B1(KEYINPUT57), .B2(new_n883), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n362), .A4(new_n841), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n875), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n890), .ZN(G1345gat));
  AOI21_X1  g690(.A(G155gat), .B1(new_n867), .B2(new_n386), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n852), .A2(new_n855), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n385), .A2(new_n430), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n867), .B2(new_n696), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n414), .A2(new_n431), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n893), .B2(new_n897), .ZN(G1347gat));
  AOI21_X1  g697(.A(new_n675), .B1(new_n819), .B2(new_n820), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n671), .A2(new_n565), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT119), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n528), .A3(new_n293), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n487), .A2(KEYINPUT120), .A3(new_n678), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n487), .B2(new_n678), .ZN(new_n905));
  NOR4_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n595), .A4(new_n687), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n853), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n293), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n528), .B2(new_n908), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n902), .B2(new_n362), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n363), .A2(new_n527), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n907), .B2(new_n911), .ZN(G1349gat));
  AOI21_X1  g711(.A(new_n386), .B1(new_n814), .B2(new_n817), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n385), .A2(new_n696), .A3(new_n293), .A4(new_n362), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n386), .B(new_n906), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n386), .A4(new_n906), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n540), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n385), .A2(new_n524), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n901), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n919), .A2(new_n925), .A3(new_n921), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n919), .B2(new_n921), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(KEYINPUT60), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT123), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n923), .B1(new_n929), .B2(new_n931), .ZN(G1350gat));
  INV_X1    g731(.A(G190gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n907), .B2(new_n696), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT61), .Z(new_n935));
  NAND3_X1  g734(.A1(new_n902), .A2(new_n933), .A3(new_n696), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1351gat));
  NOR3_X1   g736(.A1(new_n904), .A2(new_n905), .A3(new_n633), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  NAND3_X1  g738(.A1(new_n888), .A2(new_n293), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(G197gat), .A3(new_n942), .ZN(new_n943));
  AND4_X1   g742(.A1(new_n678), .A2(new_n899), .A3(new_n595), .A4(new_n634), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n489), .A3(new_n293), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(new_n362), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT62), .Z(new_n950));
  AND3_X1   g749(.A1(new_n888), .A2(new_n362), .A3(new_n939), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n948), .B2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n944), .A2(new_n376), .A3(new_n386), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n888), .A2(new_n386), .A3(new_n939), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n944), .A2(new_n492), .A3(new_n696), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n888), .A2(new_n696), .A3(new_n939), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n492), .ZN(G1355gat));
endmodule


