//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT78), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT79), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n195), .A2(new_n191), .A3(KEYINPUT79), .A4(G104), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n197), .A2(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n191), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AND4_X1   g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .A4(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n210), .A2(G128), .B1(new_n206), .B2(new_n208), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G128), .A3(new_n210), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n199), .A3(new_n202), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  INV_X1    g037(.A(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G137), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n224), .B2(G137), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n223), .A3(new_n228), .A4(new_n225), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n223), .A3(new_n225), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n230), .A2(new_n223), .A3(KEYINPUT66), .A4(new_n225), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(G131), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n221), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT12), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n221), .A2(KEYINPUT12), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n201), .B1(KEYINPUT3), .B2(new_n192), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n194), .B1(new_n248), .B2(new_n196), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n193), .A2(new_n196), .A3(new_n198), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n252), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n199), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n251), .A2(G101), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n260), .B2(new_n217), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n215), .A2(KEYINPUT64), .A3(new_n258), .A4(new_n259), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n217), .A2(KEYINPUT0), .A3(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n220), .A2(KEYINPUT10), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n199), .A2(new_n202), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n219), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n254), .A2(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n234), .A2(KEYINPUT82), .A3(new_n239), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n245), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(G227), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n277), .B(new_n279), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n270), .B2(new_n274), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n254), .A2(new_n265), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n269), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n240), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n276), .A2(new_n281), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G469), .B1(new_n287), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n221), .A2(KEYINPUT12), .A3(new_n240), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT12), .B1(new_n221), .B2(new_n240), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n243), .A2(KEYINPUT83), .A3(new_n244), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n282), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n280), .B1(new_n286), .B2(new_n275), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n289), .B(new_n291), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n190), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT2), .A2(G113), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT2), .A2(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G119), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(KEYINPUT68), .A3(new_n304), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  INV_X1    g127(.A(new_n304), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n315), .A3(new_n310), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(new_n316), .B2(KEYINPUT69), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n312), .A2(new_n315), .A3(new_n318), .A4(new_n310), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n256), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n254), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n305), .A2(new_n310), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT5), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n323), .B(G113), .C1(KEYINPUT5), .C2(new_n307), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n267), .A2(KEYINPUT84), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n324), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n203), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(G110), .B(G122), .Z(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n333));
  INV_X1    g147(.A(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(new_n334), .A3(new_n329), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT6), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n264), .A2(G125), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(G125), .B2(new_n219), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n278), .A2(G224), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(KEYINPUT6), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n334), .B1(new_n321), .B2(new_n329), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT85), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n336), .B(new_n340), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n267), .B(new_n327), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n331), .B(KEYINPUT8), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n339), .A2(KEYINPUT86), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n338), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n338), .B2(new_n352), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n355), .B2(new_n335), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n346), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n347), .B1(new_n346), .B2(new_n356), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n300), .B(new_n301), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G113), .B(G122), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n197), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  INV_X1    g178(.A(G125), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G140), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n364), .B2(new_n366), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT19), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n366), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n365), .A2(G140), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n363), .A2(G125), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT87), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n379), .B2(KEYINPUT19), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n205), .B(new_n372), .C1(new_n380), .C2(new_n371), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n384), .A3(G146), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G237), .A2(G953), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n388));
  AOI21_X1  g202(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n389));
  OAI21_X1  g203(.A(G131), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n228), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n386), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT18), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n205), .B1(new_n377), .B2(new_n378), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n373), .A2(G146), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n397), .B1(new_n390), .B2(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n362), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  AOI21_X1  g217(.A(G146), .B1(new_n382), .B2(new_n384), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n386), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT17), .B(G131), .C1(new_n388), .C2(new_n389), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n382), .A2(new_n384), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n205), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n406), .A3(new_n403), .A4(new_n385), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n393), .A2(new_n390), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n362), .B(new_n401), .C1(new_n407), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n406), .A3(new_n385), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT89), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n412), .A3(new_n410), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(KEYINPUT90), .A3(new_n362), .A4(new_n401), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n402), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT20), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n416), .A2(new_n420), .ZN(new_n427));
  INV_X1    g241(.A(new_n402), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n422), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NOR4_X1   g246(.A1(new_n421), .A2(KEYINPUT91), .A3(KEYINPUT20), .A4(new_n423), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G475), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n419), .A2(new_n401), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n427), .B1(new_n362), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G902), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT73), .B(G217), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n187), .A2(new_n278), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(KEYINPUT92), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(KEYINPUT92), .ZN(new_n447));
  OAI21_X1  g261(.A(G116), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n445), .A2(G116), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n444), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n444), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n191), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n449), .B(KEYINPUT14), .Z(new_n455));
  INV_X1    g269(.A(new_n448), .ZN(new_n456));
  OAI21_X1  g270(.A(G107), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(G128), .B(G143), .Z(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(G134), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n207), .A2(G128), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n224), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n458), .ZN(new_n464));
  INV_X1    g278(.A(new_n453), .ZN(new_n465));
  OAI21_X1  g279(.A(G107), .B1(new_n465), .B2(new_n451), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n466), .B2(new_n454), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n443), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n454), .ZN(new_n469));
  INV_X1    g283(.A(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n472));
  INV_X1    g286(.A(new_n443), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n291), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G952), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  INV_X1    g295(.A(G234), .ZN(new_n482));
  INV_X1    g296(.A(G237), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT94), .Z(new_n485));
  XOR2_X1   g299(.A(KEYINPUT21), .B(G898), .Z(new_n486));
  OAI211_X1 g300(.A(new_n290), .B(G953), .C1(new_n482), .C2(new_n483), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n475), .B(new_n291), .C1(KEYINPUT15), .C2(new_n477), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n479), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n435), .A2(new_n441), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n317), .A2(new_n319), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n264), .B1(new_n234), .B2(new_n239), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n222), .A2(G134), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n228), .B1(new_n495), .B2(new_n225), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n216), .B2(new_n218), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n234), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n234), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n234), .B2(new_n497), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n493), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n492), .B(new_n499), .C1(new_n503), .C2(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n387), .A2(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n194), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n506), .B(new_n507), .Z(new_n508));
  INV_X1    g322(.A(new_n492), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n494), .A2(new_n498), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g325(.A1(KEYINPUT70), .A2(KEYINPUT31), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n494), .A2(new_n509), .A3(KEYINPUT28), .A4(new_n498), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n516), .C1(new_n509), .C2(new_n503), .ZN(new_n517));
  INV_X1    g331(.A(new_n508), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n504), .A2(new_n508), .A3(new_n510), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n517), .B2(new_n518), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n508), .B1(new_n504), .B2(new_n510), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n291), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n498), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n492), .B1(new_n532), .B2(new_n493), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n510), .A2(new_n533), .A3(KEYINPUT71), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n492), .C1(new_n532), .C2(new_n493), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(KEYINPUT28), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n538), .A2(new_n528), .A3(new_n518), .ZN(new_n539));
  OAI21_X1  g353(.A(G472), .B1(new_n531), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n526), .A2(new_n527), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n442), .B1(new_n290), .B2(new_n482), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT74), .Z(new_n543));
  XOR2_X1   g357(.A(G119), .B(G128), .Z(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT24), .B(G110), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n306), .B2(G128), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT75), .B1(new_n306), .B2(G128), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n546), .B1(new_n550), .B2(G110), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n386), .A2(new_n400), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n544), .A2(new_n545), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n550), .B2(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n409), .A2(new_n385), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n553), .A2(new_n557), .A3(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT25), .B1(new_n566), .B2(new_n291), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n553), .A2(new_n557), .A3(new_n562), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n562), .B1(new_n553), .B2(new_n557), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT25), .B(new_n291), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n543), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n543), .A2(G902), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT77), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n566), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n360), .A2(new_n491), .A3(new_n541), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  INV_X1    g394(.A(new_n301), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n346), .A2(new_n356), .ZN(new_n582));
  INV_X1    g396(.A(new_n347), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n346), .A2(new_n347), .A3(new_n356), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n421), .A2(KEYINPUT20), .A3(new_n423), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n425), .B2(new_n424), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n441), .B1(new_n588), .B2(new_n433), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n476), .A2(G478), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n475), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n468), .A2(new_n474), .A3(KEYINPUT33), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n291), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n590), .B1(new_n594), .B2(G478), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n586), .A2(new_n589), .A3(new_n488), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n522), .A2(new_n291), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  INV_X1    g412(.A(new_n190), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n572), .A2(new_n576), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n299), .B2(new_n288), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n601), .A3(new_n524), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  AOI21_X1  g419(.A(new_n440), .B1(new_n431), .B2(new_n424), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n479), .A2(new_n489), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(KEYINPUT95), .A3(new_n488), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n431), .A2(new_n424), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n441), .A2(new_n609), .A3(new_n488), .A4(new_n607), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n586), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n608), .A2(new_n612), .A3(new_n586), .A4(KEYINPUT96), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n602), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n191), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  INV_X1    g434(.A(new_n524), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n522), .B2(new_n291), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n558), .B(new_n625), .Z(new_n626));
  OR2_X1    g440(.A1(new_n626), .A2(new_n574), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n572), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n360), .A2(new_n491), .A3(new_n624), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  INV_X1    g445(.A(new_n628), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n359), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n485), .B1(G900), .B2(new_n487), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n606), .A2(new_n607), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n541), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  AOI21_X1  g451(.A(new_n440), .B1(new_n432), .B2(new_n434), .ZN(new_n638));
  INV_X1    g452(.A(new_n607), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(G472), .A2(G902), .ZN(new_n641));
  INV_X1    g455(.A(new_n511), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n534), .A2(new_n518), .A3(new_n536), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(G472), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(KEYINPUT98), .B(new_n641), .C1(new_n642), .C2(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n526), .A2(new_n649), .A3(new_n527), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n584), .A2(new_n585), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n634), .B(KEYINPUT39), .Z(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n300), .A2(new_n655), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n581), .B(new_n628), .C1(new_n656), .C2(KEYINPUT40), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n651), .A2(new_n653), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND3_X1  g474(.A1(new_n589), .A2(new_n595), .A3(new_n634), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n633), .A2(new_n662), .A3(new_n541), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT99), .B(G146), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G48));
  NAND2_X1  g479(.A1(new_n286), .A2(new_n275), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n281), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n282), .A2(new_n295), .A3(new_n296), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n291), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n289), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n291), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n599), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n541), .A2(new_n677), .A3(new_n578), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n596), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT41), .B(G113), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT101), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n679), .B(new_n681), .ZN(G15));
  NAND2_X1  g496(.A1(new_n615), .A2(new_n616), .ZN(new_n683));
  INV_X1    g497(.A(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  OAI21_X1  g500(.A(new_n301), .B1(new_n357), .B2(new_n358), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n676), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n491), .A3(new_n541), .A4(new_n628), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n538), .A2(new_n518), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n521), .A3(new_n513), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n523), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n623), .A3(new_n577), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n488), .B(new_n301), .C1(new_n357), .C2(new_n358), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n695), .A2(new_n697), .A3(new_n640), .A4(new_n677), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NOR3_X1   g513(.A1(new_n694), .A2(new_n623), .A3(new_n632), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n662), .A2(new_n688), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n301), .A2(new_n300), .A3(new_n584), .A4(new_n585), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n541), .A3(new_n578), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n705), .B2(new_n661), .ZN(new_n706));
  INV_X1    g520(.A(new_n527), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT32), .B1(new_n522), .B2(new_n523), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n577), .B1(new_n709), .B2(new_n540), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n662), .A4(new_n704), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G131), .ZN(G33));
  AND4_X1   g527(.A1(new_n541), .A2(new_n704), .A3(new_n578), .A4(new_n635), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n224), .ZN(G36));
  NAND2_X1  g529(.A1(new_n638), .A2(new_n595), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n628), .C1(new_n621), .C2(new_n623), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n287), .A2(KEYINPUT45), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT102), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n287), .A2(KEYINPUT45), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(G469), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(G469), .A2(G902), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n299), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT46), .B1(new_n725), .B2(new_n726), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n599), .A3(new_n655), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n584), .A2(new_n301), .A3(new_n585), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT103), .Z(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G137), .ZN(G39));
  NOR4_X1   g550(.A1(new_n661), .A2(new_n541), .A3(new_n578), .A4(new_n732), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n730), .A2(new_n599), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n730), .B2(new_n599), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  INV_X1    g557(.A(new_n485), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n718), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(new_n695), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n653), .A2(new_n301), .A3(new_n676), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT50), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n732), .A2(new_n676), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n700), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n650), .A2(new_n485), .A3(new_n577), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n589), .A2(new_n595), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(KEYINPUT112), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n741), .ZN(new_n757));
  INV_X1    g571(.A(new_n675), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n674), .B1(new_n669), .B2(new_n291), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n190), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n739), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n763));
  INV_X1    g577(.A(new_n746), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n733), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n756), .A2(KEYINPUT51), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n745), .A2(new_n710), .A3(new_n750), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT114), .Z(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT48), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n746), .A2(new_n688), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n589), .A2(new_n595), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n752), .A2(new_n775), .A3(new_n750), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(new_n481), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n772), .A2(KEYINPUT48), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n755), .B(new_n749), .C1(new_n765), .C2(new_n762), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n781));
  OAI211_X1 g595(.A(new_n770), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n579), .B(new_n629), .C1(new_n596), .C2(new_n678), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n602), .A2(new_n696), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n441), .B(new_n607), .C1(new_n588), .C2(new_n433), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT106), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n435), .A2(new_n788), .A3(new_n441), .A4(new_n607), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n689), .A3(new_n698), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT105), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n602), .B1(new_n596), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n775), .A2(new_n697), .A3(KEYINPUT105), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n683), .A2(new_n684), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n714), .B1(new_n706), .B2(new_n711), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n606), .A2(new_n639), .A3(new_n634), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n632), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n801), .A2(new_n541), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n598), .A2(new_n628), .A3(new_n693), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n661), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n704), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n793), .A2(new_n797), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n541), .A2(new_n586), .A3(new_n300), .A4(new_n628), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n808), .A2(new_n635), .B1(new_n805), .B2(new_n688), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n632), .A2(new_n634), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n360), .A2(new_n650), .A3(new_n640), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n810), .A3(new_n663), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n663), .A2(new_n636), .A3(new_n701), .A4(new_n812), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n783), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n793), .A2(new_n797), .A3(new_n798), .A4(new_n806), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n813), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT53), .A4(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(KEYINPUT108), .B(new_n783), .C1(new_n807), .C2(new_n816), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n807), .A2(new_n816), .A3(new_n783), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n828), .B(new_n830), .C1(new_n831), .C2(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT110), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n827), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n782), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n480), .A2(new_n278), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT115), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n760), .B(KEYINPUT49), .Z(new_n840));
  OR2_X1    g654(.A1(new_n600), .A2(new_n581), .ZN(new_n841));
  OR4_X1    g655(.A1(new_n650), .A2(new_n840), .A3(new_n716), .A4(new_n841), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n837), .A2(new_n839), .B1(new_n653), .B2(new_n842), .ZN(G75));
  OAI21_X1  g657(.A(new_n830), .B1(new_n831), .B2(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n290), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n583), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n336), .B1(new_n343), .B2(new_n345), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n340), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT55), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n847), .B2(new_n848), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n278), .A2(G952), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(G51));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  INV_X1    g671(.A(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n832), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n726), .B(KEYINPUT57), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n669), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n845), .A2(new_n725), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n857), .B(new_n858), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n862), .B2(new_n669), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT117), .B1(new_n866), .B2(new_n854), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n846), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n869), .A2(new_n421), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n421), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n870), .A2(new_n871), .A3(new_n854), .ZN(G60));
  NAND2_X1  g686(.A1(G478), .A2(G902), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT59), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n834), .A2(new_n836), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n592), .A2(new_n593), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n876), .A2(KEYINPUT118), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT118), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  INV_X1    g693(.A(new_n855), .ZN(new_n880));
  INV_X1    g694(.A(new_n860), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n592), .A2(new_n593), .A3(new_n875), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT60), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n626), .B(KEYINPUT119), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n844), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n844), .A2(new_n887), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n880), .B(new_n889), .C1(new_n890), .C2(new_n566), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(KEYINPUT120), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(KEYINPUT120), .ZN(new_n894));
  MUX2_X1   g708(.A(new_n891), .B(new_n893), .S(new_n894), .Z(G66));
  AOI21_X1  g709(.A(new_n278), .B1(new_n486), .B2(G224), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n579), .A2(new_n629), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n679), .ZN(new_n899));
  INV_X1    g713(.A(new_n792), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n797), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n902), .B2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n849), .B1(G898), .B2(new_n278), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(G69));
  AOI21_X1  g719(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n499), .B1(new_n503), .B2(KEYINPUT30), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n372), .B1(new_n380), .B2(new_n371), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n809), .A2(new_n663), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n659), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n735), .A2(new_n742), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n732), .A2(new_n656), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n710), .B(new_n921), .C1(new_n790), .C2(new_n775), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n909), .B1(new_n923), .B2(new_n278), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G900), .A2(G953), .ZN(new_n928));
  INV_X1    g742(.A(new_n731), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(new_n586), .A3(new_n640), .A4(new_n710), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n798), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n920), .A2(new_n931), .A3(new_n912), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n909), .B(new_n928), .C1(new_n932), .C2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n924), .B2(new_n925), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n906), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n924), .A2(new_n925), .ZN(new_n936));
  INV_X1    g750(.A(new_n906), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n926), .A4(new_n933), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(G72));
  XNOR2_X1  g753(.A(new_n641), .B(KEYINPUT63), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n923), .B2(new_n901), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n504), .A2(new_n510), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n508), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n941), .B1(new_n932), .B2(new_n901), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n943), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n518), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n858), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n530), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n940), .B1(new_n952), .B2(new_n511), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n826), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(G57));
endmodule


