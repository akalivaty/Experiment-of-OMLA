//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT71), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n468), .A3(G125), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2105), .C1(new_n476), .C2(new_n474), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n478), .B2(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n467), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n469), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G136), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AND4_X1   g067(.A1(G2105), .A2(new_n463), .A3(new_n466), .A4(new_n468), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT72), .B1(new_n493), .B2(G126), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n482), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n472), .A2(new_n468), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND4_X1   g079(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n500), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n500), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n498), .A2(new_n510), .ZN(G164));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n514), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n517), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(new_n525), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT76), .B(G89), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n522), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n514), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n531), .A2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n534), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI221_X1 g127(.A(new_n550), .B1(new_n522), .B2(new_n551), .C1(new_n552), .C2(new_n525), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n514), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n525), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n572), .A2(G53), .A3(G543), .A4(new_n566), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n565), .B1(new_n574), .B2(KEYINPUT78), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n569), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G166), .ZN(G303));
  OAI21_X1  g154(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n580), .B1(new_n522), .B2(new_n581), .C1(new_n582), .C2(new_n525), .ZN(G288));
  AND2_X1   g158(.A1(new_n514), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT79), .Z(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n525), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT80), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n531), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n534), .A2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n516), .C2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n525), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n516), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n534), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n575), .A2(new_n577), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n553), .A2(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n606), .A2(G559), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n616), .B1(new_n618), .B2(G868), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g195(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n482), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n487), .B2(G135), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT84), .Z(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n442), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(KEYINPUT17), .ZN(new_n660));
  OAI22_X1  g235(.A1(new_n659), .A2(KEYINPUT86), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(KEYINPUT86), .B2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT87), .Z(new_n663));
  INV_X1    g238(.A(new_n653), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n655), .A2(new_n664), .A3(new_n657), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n655), .A2(new_n653), .A3(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT89), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n681), .A3(new_n678), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT90), .Z(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n487), .A2(G139), .ZN(new_n694));
  NAND2_X1  g269(.A1(G103), .A2(G2104), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G2105), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(KEYINPUT25), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n695), .A2(new_n698), .A3(G2105), .ZN(new_n699));
  INV_X1    g274(.A(G127), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n503), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G115), .B2(G2104), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n694), .B1(new_n697), .B2(new_n699), .C1(new_n702), .C2(new_n467), .ZN(new_n703));
  MUX2_X1   g278(.A(G33), .B(new_n703), .S(G29), .Z(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G2072), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(G2072), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT31), .B(G11), .ZN(new_n707));
  INV_X1    g282(.A(G28), .ZN(new_n708));
  AOI21_X1  g283(.A(G29), .B1(new_n708), .B2(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(KEYINPUT30), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n630), .B2(G29), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n705), .A2(new_n706), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G21), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G168), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G1966), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n487), .A2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n493), .A2(G129), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT26), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n461), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n719), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n718), .B2(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n716), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(G160), .A2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(G29), .B2(new_n740), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n736), .A2(G1961), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n715), .A2(new_n732), .A3(new_n734), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n720), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n720), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT99), .B(G2078), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n736), .A2(G1961), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n741), .A2(new_n737), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n743), .A2(new_n747), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n607), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G4), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n720), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n487), .A2(G140), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(G116), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n493), .B2(G128), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(new_n720), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n757), .A2(new_n758), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n716), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n554), .B2(new_n716), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1341), .Z(new_n775));
  NAND4_X1  g350(.A1(new_n759), .A2(new_n771), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n716), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1956), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n720), .A2(G35), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n720), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2090), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n776), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n754), .A2(new_n755), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n716), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(G288), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n716), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n716), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n716), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n792), .B1(G1971), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n591), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n794), .A2(G1971), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  MUX2_X1   g377(.A(G24), .B(G290), .S(G16), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT92), .B(G1986), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n720), .A2(G25), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n487), .A2(G131), .ZN(new_n807));
  INV_X1    g382(.A(G119), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n467), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n482), .A2(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n806), .B1(new_n813), .B2(new_n720), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT91), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n814), .B(new_n816), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n802), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n801), .A2(KEYINPUT93), .A3(KEYINPUT34), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT93), .B1(new_n801), .B2(KEYINPUT34), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n819), .B(new_n824), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n787), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n826), .ZN(G150));
  AOI22_X1  g404(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n516), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI221_X1 g408(.A(new_n831), .B1(new_n522), .B2(new_n832), .C1(new_n833), .C2(new_n525), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n606), .A2(new_n614), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n553), .A2(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n553), .A2(new_n834), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n837), .B1(new_n847), .B2(new_n849), .ZN(G145));
  INV_X1    g425(.A(new_n509), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT4), .B1(new_n508), .B2(KEYINPUT73), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n851), .A2(new_n852), .B1(new_n503), .B2(new_n502), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n854), .A2(KEYINPUT72), .A3(G126), .A4(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n495), .B1(new_n482), .B2(new_n496), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT105), .B1(new_n857), .B2(new_n492), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n859), .B(new_n491), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n853), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n768), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n813), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n493), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n467), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G142), .B2(new_n487), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n622), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n703), .B(new_n729), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n863), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G162), .B(new_n630), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G160), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n872), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT106), .B(G37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(G395));
  XNOR2_X1  g454(.A(new_n618), .B(new_n844), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n611), .A2(new_n607), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n606), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n884), .A3(new_n885), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n880), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n887), .B2(new_n880), .ZN(new_n891));
  XNOR2_X1  g466(.A(G166), .B(new_n591), .ZN(new_n892));
  XNOR2_X1  g467(.A(G290), .B(G288), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n892), .A2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n891), .B(new_n900), .Z(new_n901));
  MUX2_X1   g476(.A(new_n834), .B(new_n901), .S(G868), .Z(G295));
  MUX2_X1   g477(.A(new_n834), .B(new_n901), .S(G868), .Z(G331));
  NAND2_X1  g478(.A1(new_n843), .A2(G171), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n841), .A2(G301), .A3(new_n842), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G168), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G286), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n889), .A2(new_n886), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(new_n887), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n899), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n899), .B1(new_n909), .B2(new_n912), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n876), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n888), .A2(new_n884), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n912), .B1(new_n921), .B2(new_n910), .ZN(new_n922));
  INV_X1    g497(.A(new_n899), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n913), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n915), .C2(new_n916), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n924), .A2(KEYINPUT111), .A3(new_n925), .A4(new_n913), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n919), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n925), .B1(new_n915), .B2(new_n916), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(KEYINPUT43), .A3(new_n913), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n498), .A2(new_n859), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n491), .B1(new_n855), .B2(new_n856), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n510), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n478), .A2(new_n480), .ZN(new_n945));
  INV_X1    g520(.A(new_n471), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(G40), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n768), .B(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT112), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(new_n729), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n948), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n955), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT47), .Z(new_n958));
  OR3_X1    g533(.A1(new_n955), .A2(G1986), .A3(G290), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n729), .B(G1996), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n950), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n812), .A2(new_n816), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n812), .A2(new_n816), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n961), .B(new_n962), .C1(new_n967), .C2(new_n948), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n965), .B(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n768), .A2(new_n770), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n955), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n958), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n590), .B(G1981), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT49), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  INV_X1    g554(.A(G40), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(new_n471), .C1(new_n478), .C2(new_n480), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n861), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n977), .A2(new_n978), .A3(G8), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n789), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(G1981), .B2(new_n590), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(G8), .A3(new_n982), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n528), .A2(G8), .A3(new_n529), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n939), .A2(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n861), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n979), .B1(new_n498), .B2(new_n510), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n947), .B1(new_n993), .B2(new_n939), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n861), .A2(new_n997), .A3(new_n979), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n947), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n995), .A2(new_n996), .B1(new_n1000), .B2(G2090), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n995), .A2(new_n996), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n990), .B(G8), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G288), .A2(new_n984), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n982), .A2(G8), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n984), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n982), .A2(G8), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n983), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n987), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n861), .B2(new_n979), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  INV_X1    g588(.A(new_n991), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n1013), .B(new_n1014), .C1(new_n853), .C2(new_n941), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n853), .B2(new_n941), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n981), .B1(new_n1016), .B2(KEYINPUT116), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT117), .B(G2084), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n1018), .A2(G1966), .B1(new_n1000), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(G8), .A3(G168), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n988), .B(KEYINPUT55), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1010), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(new_n1003), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n981), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n861), .A2(new_n979), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(KEYINPUT50), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n995), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1003), .A2(new_n1036), .A3(new_n1028), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1023), .B1(new_n1037), .B2(new_n1022), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1011), .B1(new_n1029), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1017), .A2(new_n1015), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1040), .B2(new_n944), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n998), .A2(new_n999), .A3(new_n1019), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1043), .B(new_n1044), .C1(new_n1035), .C2(G168), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(KEYINPUT51), .ZN(new_n1047));
  OAI211_X1 g622(.A(G8), .B(new_n1047), .C1(new_n1021), .C2(G286), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1021), .A2(G8), .A3(G286), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1003), .A2(new_n1036), .A3(new_n1028), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT126), .ZN(new_n1053));
  INV_X1    g628(.A(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n992), .A2(new_n994), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1961), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1000), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1056), .A2(G2078), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1040), .A2(new_n944), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT62), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1037), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1053), .B1(new_n1072), .B2(new_n1051), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1039), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n992), .A2(new_n994), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1032), .A2(G1956), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n575), .B2(new_n577), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n565), .A2(KEYINPUT118), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n569), .B2(new_n573), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n565), .A2(KEYINPUT118), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT119), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1081), .A2(new_n1086), .A3(KEYINPUT119), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1078), .A2(new_n1079), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1032), .A2(G1956), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1089), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1087), .A3(new_n1092), .A4(new_n1077), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n982), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n758), .A2(new_n1000), .B1(new_n1095), .B2(new_n770), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n606), .B1(new_n1096), .B2(KEYINPUT60), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n992), .A2(new_n994), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  OAI22_X1  g676(.A1(G1996), .A2(new_n1100), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n554), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1093), .A2(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1092), .A2(new_n1110), .A3(new_n1087), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(new_n1079), .C2(new_n1078), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n606), .B2(new_n1096), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1099), .A2(new_n1114), .B1(new_n1093), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1118));
  AOI21_X1  g693(.A(G171), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  AND4_X1   g696(.A1(G40), .A2(new_n946), .A3(new_n477), .A4(new_n1060), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n992), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1123), .B2(new_n1012), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n944), .A2(KEYINPUT123), .A3(new_n992), .A4(new_n1122), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1059), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1057), .ZN(new_n1127));
  OAI21_X1  g702(.A(G171), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1052), .A2(new_n1069), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1119), .A2(new_n1059), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1065), .A2(new_n1066), .A3(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1132), .A2(KEYINPUT124), .A3(new_n1117), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT124), .B1(new_n1132), .B2(new_n1117), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1116), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1130), .B(KEYINPUT125), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1074), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n967), .A2(new_n948), .ZN(new_n1140));
  XOR2_X1   g715(.A(G290), .B(G1986), .Z(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n955), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT113), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n973), .B1(new_n1139), .B2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g719(.A1(new_n458), .A2(new_n692), .A3(new_n651), .A4(new_n670), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n931), .A2(new_n877), .A3(new_n1146), .ZN(G225));
  INV_X1    g721(.A(G225), .ZN(G308));
endmodule


