//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(G244), .Z(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n211), .B1(new_n214), .B2(new_n216), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT12), .ZN(new_n245));
  OR2_X1    g0045(.A1(KEYINPUT67), .A2(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT67), .A2(G1), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n246), .A2(G13), .A3(G20), .A4(new_n247), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n245), .B1(new_n248), .B2(G68), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT67), .A2(G1), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT67), .A2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n253), .A2(KEYINPUT12), .A3(G13), .A4(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n212), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n246), .A2(new_n247), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(G68), .C1(new_n259), .C2(new_n252), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n249), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT11), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n254), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n252), .A2(G33), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n266), .B(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n257), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n270), .B2(new_n257), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n264), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n274), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n277));
  AND4_X1   g0077(.A1(new_n262), .A2(new_n263), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(G226), .A4(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT70), .A3(G226), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n283), .A2(new_n285), .A3(G232), .A4(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G97), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n282), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G41), .A2(G45), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G1), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n282), .A2(new_n299), .A3(G274), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n282), .B1(new_n259), .B2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(G238), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT13), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n300), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n250), .A2(new_n251), .ZN(new_n307));
  INV_X1    g0107(.A(new_n298), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n305), .B1(new_n309), .B2(G238), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n295), .B1(new_n289), .B2(new_n291), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n282), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n304), .A2(new_n313), .A3(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n315), .B1(new_n314), .B2(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n279), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n300), .B1(new_n301), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n290), .A2(G222), .A3(new_n286), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n283), .A2(new_n285), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G77), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n290), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n324), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n306), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT68), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(new_n300), .C1(new_n301), .C2(new_n321), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n323), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n248), .A2(G50), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n253), .A2(new_n257), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(G50), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT8), .B(G58), .Z(new_n339));
  INV_X1    g0139(.A(KEYINPUT69), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  INV_X1    g0143(.A(new_n269), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n338), .B1(new_n347), .B2(new_n258), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n323), .A2(new_n330), .A3(new_n349), .A4(new_n332), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n335), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(KEYINPUT9), .B(new_n338), .C1(new_n347), .C2(new_n258), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  INV_X1    g0153(.A(new_n338), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n258), .B1(new_n345), .B2(new_n346), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT10), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n333), .A2(G200), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n323), .A2(new_n330), .A3(G190), .A4(new_n332), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n352), .A2(new_n356), .A3(new_n360), .ZN(new_n362));
  INV_X1    g0162(.A(new_n359), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT10), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n351), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n217), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n300), .B1(new_n301), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n290), .A2(G232), .A3(new_n286), .ZN(new_n368));
  INV_X1    g0168(.A(G107), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n369), .B2(new_n290), .C1(new_n327), .C2(new_n302), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n306), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(G169), .ZN(new_n372));
  INV_X1    g0172(.A(new_n265), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n342), .A2(new_n373), .B1(new_n252), .B2(new_n268), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n269), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n257), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n337), .A2(G77), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(G77), .C2(new_n248), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n371), .A2(new_n349), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n372), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n371), .B2(G190), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n371), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n314), .A2(G200), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n304), .A2(new_n313), .A3(G190), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n278), .A3(new_n387), .ZN(new_n388));
  AND4_X1   g0188(.A1(new_n320), .A2(new_n365), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n328), .A2(new_n286), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n321), .A2(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n283), .A2(new_n390), .A3(new_n285), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n392), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT74), .B1(new_n392), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n306), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT75), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n306), .C1(new_n394), .C2(new_n395), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n300), .B1(new_n301), .B2(new_n233), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(G190), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n395), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n392), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n282), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n383), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G58), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n254), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n409), .A2(new_n201), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n290), .B2(G20), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n252), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n254), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(KEYINPUT73), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(new_n254), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT16), .B(new_n411), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(new_n411), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n422), .A3(new_n257), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n341), .A2(new_n343), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n257), .B2(new_n253), .ZN(new_n425));
  INV_X1    g0225(.A(new_n248), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n424), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n407), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n407), .A2(new_n423), .A3(KEYINPUT78), .A4(new_n427), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n434), .B2(KEYINPUT17), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT77), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n400), .A2(G179), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n397), .A2(new_n399), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n334), .B1(new_n405), .B2(new_n400), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n423), .A2(new_n427), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n443), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT18), .A4(new_n444), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n436), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT77), .B1(new_n445), .B2(new_n446), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n389), .B(new_n435), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n438), .A2(new_n443), .A3(new_n439), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n443), .B1(new_n438), .B2(new_n439), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT18), .B1(new_n456), .B2(new_n442), .ZN(new_n457));
  INV_X1    g0257(.A(new_n448), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT77), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(KEYINPUT79), .A3(new_n435), .A4(new_n389), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT81), .B1(new_n464), .B2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n281), .A3(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n246), .A2(G45), .A3(new_n247), .ZN(new_n471));
  OAI211_X1 g0271(.A(G270), .B(new_n282), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n283), .A2(new_n285), .A3(G264), .A4(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n283), .A2(new_n285), .A3(G257), .A4(new_n286), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT85), .B(G303), .Z(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n290), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n306), .ZN(new_n478));
  INV_X1    g0278(.A(G274), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n306), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n465), .A2(new_n467), .B1(new_n464), .B2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n250), .A2(new_n251), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(G270), .A4(new_n282), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n473), .A2(new_n478), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n487), .A2(new_n484), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(G190), .A3(new_n478), .A4(new_n473), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n280), .B2(G97), .ZN(new_n492));
  NAND3_X1  g0292(.A1(KEYINPUT80), .A2(G33), .A3(G283), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT80), .B1(G33), .B2(G283), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n256), .A2(new_n212), .B1(G20), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n496), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT20), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n246), .A2(G33), .A3(new_n247), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n248), .A2(new_n258), .A3(new_n501), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n499), .A2(new_n500), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT86), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n426), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT86), .B1(new_n248), .B2(G116), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n489), .A2(new_n491), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n349), .B1(new_n477), .B2(new_n306), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n503), .B2(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n473), .A2(new_n484), .A3(new_n487), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n487), .A2(new_n484), .ZN(new_n515));
  INV_X1    g0315(.A(new_n478), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n306), .B1(new_n481), .B2(new_n483), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n486), .B1(new_n517), .B2(G270), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G169), .B1(new_n503), .B2(new_n507), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT21), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  INV_X1    g0322(.A(new_n500), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n496), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n524));
  INV_X1    g0324(.A(new_n502), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n505), .A2(new_n506), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n334), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n522), .B1(new_n528), .B2(new_n488), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n509), .B(new_n514), .C1(new_n521), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n483), .A2(new_n468), .A3(new_n469), .ZN(new_n532));
  AOI22_X1  g0332(.A1(G257), .A2(new_n517), .B1(new_n532), .B2(new_n480), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(new_n286), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n494), .A2(new_n495), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n306), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n533), .A2(new_n534), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n534), .B1(new_n533), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(G190), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n369), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n369), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n205), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(KEYINPUT6), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n413), .A2(new_n414), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n258), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n426), .A2(new_n547), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n547), .B2(new_n502), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(new_n282), .C1(new_n470), .C2(new_n471), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n558), .A2(new_n559), .A3(new_n484), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n558), .B2(new_n484), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n542), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G200), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n545), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n541), .A2(new_n306), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n558), .A2(new_n484), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT83), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n533), .A2(new_n534), .A3(new_n542), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n334), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n349), .B(new_n542), .C1(new_n560), .C2(new_n561), .ZN(new_n570));
  INV_X1    g0370(.A(new_n557), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n283), .A2(new_n285), .A3(new_n252), .A4(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT88), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n290), .A2(new_n577), .A3(new_n252), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n252), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n369), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n344), .A2(G116), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n574), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n580), .B1(new_n576), .B2(new_n578), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n574), .B(new_n588), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n257), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n248), .A2(G107), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n595), .A2(KEYINPUT25), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(KEYINPUT25), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(G107), .B2(new_n525), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n517), .A2(G264), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G294), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n283), .A2(new_n285), .A3(G250), .A4(new_n286), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n306), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n604), .A3(new_n484), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n383), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G190), .B2(new_n605), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n594), .A2(new_n598), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n605), .A2(G179), .ZN(new_n609));
  AOI22_X1  g0409(.A1(G264), .A2(new_n517), .B1(new_n603), .B2(new_n306), .ZN(new_n610));
  AOI21_X1  g0410(.A(G169), .B1(new_n610), .B2(new_n484), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT24), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n258), .B1(new_n614), .B2(new_n592), .ZN(new_n615));
  INV_X1    g0415(.A(new_n598), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n375), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n248), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n252), .B1(new_n294), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G87), .B2(new_n206), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n283), .A2(new_n285), .A3(new_n252), .A4(G68), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n269), .B2(new_n547), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n625), .B2(new_n257), .ZN(new_n626));
  INV_X1    g0426(.A(G87), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n502), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n290), .A2(G244), .A3(G1698), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G33), .A2(G116), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n283), .A2(new_n285), .A3(G238), .A4(new_n286), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n246), .A2(G45), .A3(new_n479), .A4(new_n247), .ZN(new_n633));
  INV_X1    g0433(.A(G250), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n306), .B1(new_n471), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n632), .A2(new_n306), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n628), .B1(G190), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n383), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n525), .A2(new_n618), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n349), .A2(new_n636), .B1(new_n626), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n306), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n282), .B(new_n633), .C1(new_n483), .C2(G250), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n334), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n637), .A2(new_n639), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n608), .A2(new_n617), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n463), .A2(new_n531), .A3(new_n573), .A4(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n635), .A2(new_n650), .A3(new_n633), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n334), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n641), .A2(new_n645), .ZN(new_n656));
  INV_X1    g0456(.A(G190), .ZN(new_n657));
  OAI221_X1 g0457(.A(new_n626), .B1(new_n627), .B2(new_n502), .C1(new_n644), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(new_n638), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n572), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT21), .B1(new_n519), .B2(new_n520), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n528), .A2(new_n522), .A3(new_n488), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n514), .ZN(new_n667));
  AOI211_X1 g0467(.A(KEYINPUT90), .B(new_n513), .C1(new_n664), .C2(new_n665), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n617), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n652), .A2(G200), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n654), .B1(new_n637), .B2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n572), .A2(new_n671), .A3(new_n564), .A4(new_n608), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n662), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n569), .A2(new_n570), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT91), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n569), .A2(new_n676), .A3(new_n570), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n571), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n675), .A2(KEYINPUT92), .A3(new_n571), .A4(new_n677), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n661), .A3(new_n681), .A4(new_n671), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n463), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n388), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n320), .B1(new_n685), .B2(new_n381), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n435), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n447), .A2(new_n448), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n361), .A2(new_n364), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n351), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(G369));
  NOR2_X1   g0493(.A1(new_n667), .A2(new_n668), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n252), .A2(G13), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n307), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n508), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n530), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n608), .A2(new_n617), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n701), .B1(new_n615), .B2(new_n616), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n617), .B2(new_n702), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n666), .A2(new_n514), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n702), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(new_n708), .ZN(new_n716));
  INV_X1    g0516(.A(new_n617), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n702), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n209), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n216), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n701), .B1(new_n673), .B2(new_n682), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n671), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n678), .B2(new_n679), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n661), .B1(new_n731), .B2(new_n681), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n617), .A2(new_n666), .A3(new_n514), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n672), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n701), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n647), .A2(new_n573), .A3(new_n531), .A4(new_n702), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n567), .A2(new_n568), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n610), .A2(new_n510), .A3(new_n636), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n512), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n743), .A2(KEYINPUT30), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT30), .B1(new_n743), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n566), .A2(KEYINPUT82), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n558), .A2(new_n559), .A3(new_n484), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n565), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n605), .A2(new_n652), .A3(new_n349), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n750), .A2(new_n519), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n742), .B1(new_n753), .B2(new_n702), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n743), .A2(new_n745), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n750), .A2(new_n751), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(KEYINPUT30), .B1(new_n756), .B2(new_n519), .ZN(new_n757));
  OAI211_X1 g0557(.A(KEYINPUT31), .B(new_n701), .C1(new_n757), .C2(new_n746), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n741), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n740), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n726), .B1(new_n762), .B2(G1), .ZN(G364));
  INV_X1    g0563(.A(G1), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n695), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n721), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n707), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n705), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n290), .A2(new_n209), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n209), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n240), .A2(new_n482), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n720), .A2(new_n290), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n216), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(new_n482), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n772), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n252), .B1(KEYINPUT93), .B2(new_n334), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(KEYINPUT93), .B2(new_n334), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n213), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n767), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n252), .A2(new_n349), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n252), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n792), .A2(new_n408), .B1(new_n794), .B2(new_n627), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n790), .A2(new_n383), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n202), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G190), .A2(G200), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n789), .A2(new_n657), .A3(G200), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n290), .B1(new_n800), .B2(new_n268), .C1(new_n254), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n793), .A2(new_n657), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n369), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n795), .A2(new_n798), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n349), .A2(new_n383), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n252), .A2(G190), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n252), .B1(new_n808), .B2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G97), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT32), .B1(new_n810), .B2(new_n811), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n805), .A2(new_n812), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G322), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n792), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G326), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n797), .A2(new_n822), .B1(new_n803), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n794), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n821), .B(new_n824), .C1(G303), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n810), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G329), .ZN(new_n828));
  INV_X1    g0628(.A(new_n800), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(G311), .ZN(new_n830));
  INV_X1    g0630(.A(new_n801), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n290), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n826), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n817), .B1(new_n819), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n788), .B1(new_n835), .B2(new_n782), .ZN(new_n836));
  INV_X1    g0636(.A(new_n785), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n705), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n769), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  OAI21_X1  g0640(.A(new_n815), .B1(new_n818), .B2(new_n792), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT95), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n325), .B1(new_n800), .B2(new_n497), .C1(new_n823), .C2(new_n801), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n803), .A2(new_n627), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G303), .B2(new_n796), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n369), .B2(new_n794), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(G311), .C2(new_n827), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n290), .B1(new_n803), .B2(new_n254), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G50), .B2(new_n825), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n408), .B2(new_n813), .C1(new_n852), .C2(new_n810), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n831), .A2(G150), .B1(new_n829), .B2(G159), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT97), .B(G143), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(new_n792), .B2(new_n855), .C1(new_n856), .C2(new_n797), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  OAI21_X1  g0658(.A(new_n849), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n782), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n781), .A2(new_n784), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(new_n767), .C1(G77), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n381), .A2(new_n701), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n701), .A2(new_n379), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n384), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n381), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n783), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n869), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n727), .B(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(new_n760), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n767), .B1(new_n872), .B2(new_n760), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  NOR2_X1   g0676(.A1(new_n278), .A2(new_n702), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n320), .A2(new_n388), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n314), .A2(G169), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT14), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n388), .A2(new_n881), .A3(new_n317), .A4(new_n316), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT99), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n877), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n869), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n759), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n741), .A2(new_n754), .A3(new_n758), .A4(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n699), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n442), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n445), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(new_n434), .ZN(new_n898));
  INV_X1    g0698(.A(new_n427), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n419), .A2(new_n257), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n411), .B1(new_n416), .B2(new_n418), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n420), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n441), .A2(new_n444), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n699), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n434), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n435), .B1(new_n449), .B2(new_n450), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n903), .A2(new_n699), .ZN(new_n908));
  AOI221_X4 g0708(.A(new_n893), .B1(new_n898), .B2(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n906), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n892), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n896), .B1(new_n435), .B2(new_n688), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n434), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT37), .B1(new_n456), .B2(new_n442), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT100), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n896), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n445), .A2(new_n428), .A3(new_n896), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT100), .B1(new_n897), .B2(new_n434), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n892), .B(KEYINPUT40), .C1(new_n909), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n916), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n889), .A2(new_n891), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n463), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n929), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n909), .B2(new_n927), .ZN(new_n935));
  INV_X1    g0735(.A(new_n908), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n461), .B2(new_n435), .ZN(new_n937));
  INV_X1    g0737(.A(new_n911), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n893), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n320), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n702), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n688), .A2(new_n895), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n939), .A2(new_n940), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n887), .A2(new_n879), .A3(new_n884), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n727), .A2(new_n871), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n865), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n691), .A2(new_n351), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n739), .B2(new_n463), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n953), .B(new_n955), .Z(new_n956));
  OAI22_X1  g0756(.A1(new_n933), .A2(new_n956), .B1(new_n307), .B2(new_n695), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n933), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n214), .A2(new_n497), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n550), .B2(KEYINPUT35), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT98), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n961), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT36), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n216), .A2(new_n268), .A3(new_n409), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n202), .A2(G68), .ZN(new_n967));
  AOI211_X1 g0767(.A(G13), .B(new_n307), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n958), .A2(new_n965), .A3(new_n968), .ZN(G367));
  OR2_X1    g0769(.A1(new_n678), .A2(new_n702), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n573), .B1(new_n557), .B2(new_n702), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n716), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT42), .Z(new_n974));
  AOI21_X1  g0774(.A(new_n617), .B1(new_n970), .B2(new_n971), .ZN(new_n975));
  INV_X1    g0775(.A(new_n572), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n702), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n701), .A2(new_n628), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n654), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n730), .B2(new_n980), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT103), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n978), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  MUX2_X1   g0786(.A(new_n978), .B(new_n984), .S(new_n986), .Z(new_n987));
  AOI21_X1  g0787(.A(new_n712), .B1(new_n971), .B2(new_n970), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT105), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n718), .A2(new_n972), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT45), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n718), .A2(new_n972), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT44), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n712), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT107), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n716), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n711), .A2(new_n715), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n707), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n761), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1000), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n762), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n721), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n994), .B1(new_n1015), .B2(new_n766), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n231), .A2(new_n775), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n786), .B1(new_n209), .B2(new_n375), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n767), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n325), .B1(new_n831), .B2(G159), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n202), .B2(new_n800), .C1(new_n810), .C2(new_n856), .ZN(new_n1021));
  INV_X1    g0821(.A(G150), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n792), .A2(new_n1022), .B1(new_n803), .B2(new_n268), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n797), .A2(new_n855), .B1(new_n408), .B2(new_n794), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n254), .B2(new_n813), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT46), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n794), .A2(new_n1027), .A3(new_n497), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT108), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n325), .B1(new_n800), .B2(new_n823), .C1(new_n818), .C2(new_n801), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n827), .B2(G317), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n792), .A2(new_n476), .B1(new_n803), .B2(new_n547), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G311), .B2(new_n796), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n814), .A2(G107), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1027), .B1(new_n794), .B2(new_n497), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT47), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1019), .B1(new_n1038), .B2(new_n782), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n983), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n837), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1016), .A2(new_n1041), .ZN(G387));
  NAND2_X1  g0842(.A1(new_n1007), .A2(new_n761), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1010), .A2(new_n721), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1007), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n711), .A2(new_n837), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n236), .A2(new_n482), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT109), .Z(new_n1048));
  NOR2_X1   g0848(.A1(new_n342), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n482), .B1(new_n254), .B2(new_n268), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n775), .B(new_n1048), .C1(new_n1050), .C2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n723), .A2(new_n771), .B1(G107), .B2(new_n209), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n786), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n767), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n290), .B1(new_n800), .B2(new_n254), .C1(new_n547), .C2(new_n803), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n827), .B2(G150), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n814), .A2(new_n618), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n825), .A2(G77), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n797), .B2(new_n811), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G50), .B2(new_n791), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n424), .A2(new_n831), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n476), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G311), .A2(new_n831), .B1(new_n1067), .B2(new_n829), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n791), .A2(G317), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n820), .C2(new_n797), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n823), .B2(new_n813), .C1(new_n818), .C2(new_n794), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT49), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n325), .B1(new_n497), .B2(new_n803), .C1(new_n810), .C2(new_n822), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1058), .B1(new_n1078), .B2(new_n782), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1045), .A2(new_n766), .B1(new_n1046), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1044), .A2(new_n1080), .ZN(G393));
  OAI21_X1  g0881(.A(new_n786), .B1(new_n547), .B2(new_n209), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n243), .A2(new_n775), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n767), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT113), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n972), .A2(new_n837), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT112), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n325), .B1(new_n800), .B2(new_n818), .C1(new_n476), .C2(new_n801), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n804), .B(new_n1088), .C1(G283), .C2(new_n825), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n497), .B2(new_n813), .C1(new_n820), .C2(new_n810), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n791), .B1(new_n796), .B2(G317), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G150), .A2(new_n796), .B1(new_n791), .B2(G159), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n290), .B1(new_n800), .B2(new_n342), .C1(new_n202), .C2(new_n801), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n844), .B(new_n1095), .C1(G68), .C2(new_n825), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n814), .A2(G77), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n810), .C2(new_n855), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1090), .A2(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1085), .B(new_n1087), .C1(new_n782), .C2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n765), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n721), .B1(new_n1008), .B2(new_n1000), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(G390));
  NAND4_X1  g0906(.A1(new_n888), .A2(new_n889), .A3(G330), .A4(new_n891), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n701), .B(new_n869), .C1(new_n673), .C2(new_n682), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n948), .B1(new_n1109), .B2(new_n864), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n935), .A2(new_n941), .B1(new_n1110), .B2(new_n943), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n893), .B1(new_n1112), .B2(new_n917), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n944), .B1(new_n1113), .B2(new_n940), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n702), .B(new_n868), .C1(new_n732), .C2(new_n736), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n865), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n948), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1110), .A2(new_n943), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n909), .A2(new_n912), .A3(new_n934), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT39), .B1(new_n1113), .B2(new_n940), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n759), .A2(new_n948), .A3(G330), .A4(new_n871), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n766), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n783), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n767), .B1(new_n424), .B2(new_n862), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT117), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n497), .A2(new_n792), .B1(new_n797), .B2(new_n823), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n254), .A2(new_n803), .B1(new_n794), .B2(new_n627), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n827), .A2(G294), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n325), .B1(new_n800), .B2(new_n547), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G107), .B2(new_n831), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1097), .A2(new_n1134), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n794), .A2(new_n1022), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n290), .B1(new_n800), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G137), .B2(new_n831), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1140), .B(new_n1143), .C1(new_n1144), .C2(new_n810), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n796), .A2(G128), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n803), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n791), .A2(G132), .B1(new_n1147), .B2(G50), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(new_n813), .C2(new_n811), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1138), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1131), .B1(new_n1150), .B2(new_n782), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1129), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1128), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT114), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n950), .A2(new_n865), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n949), .B1(new_n760), .B2(new_n869), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1107), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1115), .A2(new_n865), .A3(new_n1125), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n889), .A2(G330), .A3(new_n871), .A4(new_n891), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n949), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1156), .A2(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n660), .A2(new_n661), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n655), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n672), .B2(new_n733), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n680), .A2(new_n681), .A3(new_n671), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n661), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n728), .B1(new_n1167), .B2(new_n702), .ZN(new_n1168));
  AOI211_X1 g0968(.A(KEYINPUT29), .B(new_n701), .C1(new_n673), .C2(new_n682), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n463), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n463), .A2(new_n930), .A3(G330), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n692), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1155), .B1(new_n1162), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1158), .A2(new_n1156), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1176), .A2(new_n955), .A3(KEYINPUT114), .A4(new_n1171), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n722), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT115), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1178), .A2(new_n1181), .A3(new_n1179), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT115), .B1(new_n1127), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(KEYINPUT116), .B(new_n1180), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1127), .A2(KEYINPUT115), .A3(new_n1183), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT116), .B1(new_n1189), .B2(new_n1180), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1154), .B1(new_n1186), .B2(new_n1190), .ZN(G378));
  NAND2_X1  g0991(.A1(new_n348), .A2(new_n895), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n365), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n365), .A2(new_n1192), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n783), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n767), .B1(new_n862), .B2(G50), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n791), .A2(G128), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n794), .B2(new_n1141), .C1(new_n797), .C2(new_n1144), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n801), .A2(new_n852), .B1(new_n800), .B2(new_n856), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT119), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G150), .C2(new_n814), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n280), .B(new_n281), .C1(new_n803), .C2(new_n811), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n827), .B2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n290), .A2(G41), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n800), .B2(new_n375), .C1(new_n547), .C2(new_n801), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1062), .B1(new_n792), .B2(new_n369), .C1(new_n497), .C2(new_n797), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G283), .C2(new_n827), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n803), .A2(new_n408), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT118), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n254), .C2(new_n813), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1214), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1213), .A2(new_n1222), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1202), .B1(new_n1226), .B2(new_n782), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n939), .B2(new_n940), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n928), .B(G330), .C1(new_n1231), .C2(new_n914), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1200), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n916), .A2(new_n1199), .A3(G330), .A4(new_n928), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n953), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT121), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1233), .A2(new_n953), .A3(new_n1234), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT120), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n953), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT121), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(KEYINPUT120), .ZN(new_n1245));
  AOI211_X1 g1045(.A(KEYINPUT121), .B(new_n953), .C1(new_n1234), .C2(new_n1233), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1244), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1229), .B1(new_n1249), .B2(new_n766), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n955), .B(new_n1171), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1172), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT57), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n721), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1250), .B1(new_n1252), .B2(new_n1256), .ZN(G375));
  NAND2_X1  g1057(.A1(new_n949), .A2(new_n783), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n767), .B1(new_n862), .B2(G68), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n823), .A2(new_n792), .B1(new_n797), .B2(new_n818), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n268), .A2(new_n803), .B1(new_n794), .B2(new_n547), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n827), .A2(G303), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n325), .B1(new_n800), .B2(new_n369), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G116), .B2(new_n831), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1061), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1219), .A2(new_n290), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n814), .A2(G50), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n827), .A2(G128), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n801), .A2(new_n1141), .B1(new_n800), .B2(new_n1022), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G132), .B2(new_n796), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n791), .A2(G137), .B1(new_n825), .B2(G159), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1266), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1259), .B1(new_n1275), .B2(new_n782), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1176), .A2(new_n766), .B1(new_n1258), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1178), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1279), .B2(new_n1013), .ZN(G381));
  AND2_X1   g1080(.A1(new_n1016), .A2(new_n1041), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1153), .B1(new_n1189), .B2(new_n1180), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1044), .A2(new_n839), .A3(new_n1080), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(G375), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n700), .A2(G213), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G407), .B(G213), .C1(G375), .C2(new_n1289), .ZN(G409));
  OAI211_X1 g1090(.A(G378), .B(new_n1250), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1251), .A2(new_n1014), .A3(new_n1244), .A4(new_n1248), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1239), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n766), .B1(new_n1293), .B2(new_n1241), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT123), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1228), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(new_n1294), .B2(new_n1228), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1292), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1282), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1288), .B1(new_n1291), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1288), .A2(G2897), .ZN(new_n1302));
  XOR2_X1   g1102(.A(new_n1302), .B(KEYINPUT124), .Z(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1279), .A2(KEYINPUT60), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n722), .B1(new_n1278), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(G384), .A3(new_n1277), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1308), .B2(new_n1277), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1311), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1309), .A3(new_n1303), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(KEYINPUT125), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1318));
  OR3_X1    g1118(.A1(new_n1301), .A2(new_n1316), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n839), .B1(new_n1044), .B2(new_n1080), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G390), .A2(new_n1283), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1283), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(G387), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(KEYINPUT61), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1313), .A2(new_n1309), .ZN(new_n1328));
  AOI211_X1 g1128(.A(new_n1288), .B(new_n1328), .C1(new_n1291), .C2(new_n1300), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT63), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1301), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1319), .A2(new_n1327), .A3(new_n1330), .A4(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1301), .B2(new_n1315), .ZN(new_n1337));
  AND2_X1   g1137(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1338), .B1(new_n1329), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1332), .A2(new_n1339), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1337), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1326), .B(KEYINPUT127), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1335), .B1(new_n1343), .B2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1282), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1291), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1331), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1291), .A3(new_n1328), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1326), .ZN(G402));
endmodule


