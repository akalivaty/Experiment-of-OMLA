//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n471), .A2(KEYINPUT68), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n474), .B1(new_n483), .B2(G2105), .ZN(G160));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n485), .A2(new_n465), .A3(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n485), .B2(new_n465), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n465), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n472), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n476), .B2(new_n477), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n471), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n465), .B2(G114), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(G126), .A2(new_n490), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n502), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n515), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n528));
  INV_X1    g103(.A(new_n526), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G88), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n526), .A2(new_n517), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n536), .A2(G651), .B1(G50), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  XNOR2_X1  g115(.A(KEYINPUT75), .B(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(G76), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n529), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G51), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G63), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n523), .A2(new_n550), .B1(new_n543), .B2(new_n544), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n549), .B1(G651), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n542), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n554), .B2(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(KEYINPUT76), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n537), .A2(G52), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n527), .A2(new_n530), .ZN(new_n558));
  INV_X1    g133(.A(G90), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n556), .A2(new_n560), .ZN(G171));
  NAND2_X1  g136(.A1(new_n531), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n523), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G43), .B2(new_n537), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G53), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n547), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n547), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n523), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n577), .A2(new_n578), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n531), .A2(G91), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G299));
  OR2_X1    g159(.A1(new_n556), .A2(new_n560), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND2_X1  g162(.A1(G171), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND2_X1  g166(.A1(new_n531), .A2(G87), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n528), .A2(G74), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G49), .B2(new_n537), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n523), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G48), .B2(new_n537), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n527), .A2(G86), .A3(new_n530), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n523), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G47), .B2(new_n537), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n558), .ZN(G290));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT81), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(KEYINPUT81), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n523), .C2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n537), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n558), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT80), .B1(new_n619), .B2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n589), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n620), .B(KEYINPUT80), .S(new_n622), .Z(G321));
  XNOR2_X1  g198(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NOR2_X1   g199(.A1(G286), .A2(new_n621), .ZN(new_n625));
  XOR2_X1   g200(.A(G299), .B(KEYINPUT83), .Z(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n621), .ZN(G297));
  AOI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(new_n621), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(new_n629), .B2(G860), .ZN(G148));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n615), .A2(new_n618), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n613), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n633), .B2(G559), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n619), .A2(KEYINPUT84), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  MUX2_X1   g211(.A(new_n567), .B(new_n636), .S(G868), .Z(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n471), .A2(new_n467), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n490), .A2(G123), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n465), .A2(KEYINPUT86), .A3(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(KEYINPUT86), .B1(new_n465), .B2(G111), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G2104), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G135), .ZN(new_n651));
  OAI221_X1 g226(.A(new_n646), .B1(new_n647), .B2(new_n650), .C1(new_n651), .C2(new_n472), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n644), .A2(new_n645), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT87), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2443), .B(G2446), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(new_n670), .A3(G14), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n446), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(KEYINPUT17), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n672), .B(new_n673), .C1(new_n446), .C2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n674), .A3(new_n672), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n687), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT89), .Z(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G29), .B2(G32), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n478), .A2(G2105), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G141), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n490), .A2(G129), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n467), .A2(G105), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT26), .Z(new_n712));
  AND4_X1   g287(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n704), .B(new_n705), .S(new_n714), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  INV_X1    g291(.A(G34), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT24), .ZN(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n717), .B2(KEYINPUT24), .ZN(new_n719));
  AOI22_X1  g294(.A1(G160), .A2(G29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n715), .A2(new_n716), .B1(G2084), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G33), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n706), .A2(G139), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n726), .B(new_n727), .C1(new_n465), .C2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(new_n444), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT96), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n722), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n722), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT29), .B(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n720), .A2(G2084), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT30), .B(G28), .ZN(new_n740));
  OR2_X1    g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  NAND2_X1  g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n740), .A2(new_n722), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n652), .B2(new_n722), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n738), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NOR2_X1   g321(.A1(G171), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G5), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n745), .B1(new_n749), .B2(G1961), .C1(new_n716), .C2(new_n715), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G299), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G1956), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G1956), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n490), .A2(G128), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n465), .A2(G116), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n759));
  INV_X1    g334(.A(G140), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n757), .B1(new_n758), .B2(new_n759), .C1(new_n760), .C2(new_n472), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n722), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n722), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n722), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(new_n445), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n756), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n750), .A2(new_n755), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n746), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n568), .B2(new_n746), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1341), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n746), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n746), .ZN(new_n777));
  INV_X1    g352(.A(G1966), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n775), .B(new_n779), .C1(new_n780), .C2(new_n748), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n746), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n619), .B2(new_n746), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1348), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n734), .A2(new_n772), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n746), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n746), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n746), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n746), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  INV_X1    g373(.A(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n796), .B(new_n800), .C1(new_n795), .C2(new_n794), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n490), .A2(G119), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n465), .A2(G107), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G131), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n807), .C2(new_n472), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT90), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  INV_X1    g387(.A(G1986), .ZN(new_n813));
  INV_X1    g388(.A(G290), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n746), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n746), .B2(G24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n812), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n813), .B2(new_n816), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n802), .A2(new_n803), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n802), .A2(new_n821), .A3(new_n803), .A4(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n786), .B1(new_n820), .B2(new_n822), .ZN(G311));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(new_n786), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(G150));
  AOI22_X1  g401(.A1(new_n531), .A2(G93), .B1(G55), .B2(new_n537), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  OAI21_X1  g404(.A(G651), .B1(new_n828), .B2(KEYINPUT97), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n619), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT98), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(new_n568), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n833), .B1(new_n839), .B2(new_n841), .ZN(G145));
  XOR2_X1   g417(.A(new_n513), .B(new_n761), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n713), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n729), .ZN(new_n845));
  INV_X1    g420(.A(new_n730), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n844), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n808), .B(new_n641), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n490), .A2(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n706), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n848), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(G160), .B(KEYINPUT99), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n652), .ZN(new_n858));
  INV_X1    g433(.A(new_n854), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n845), .B(new_n859), .C1(new_n846), .C2(new_n844), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT100), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n858), .B1(new_n855), .B2(new_n860), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n837), .A2(new_n634), .A3(new_n635), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n831), .B(new_n567), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n636), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n633), .A2(new_n753), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n619), .A2(G299), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n873), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n633), .A2(new_n753), .A3(KEYINPUT101), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n878), .A3(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n633), .A2(KEYINPUT102), .A3(new_n753), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n871), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n876), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n871), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(G288), .B(G305), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n814), .B(G303), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n887), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n897), .A2(new_n884), .A3(KEYINPUT103), .A4(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G868), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n867), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n887), .A2(new_n890), .A3(new_n898), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(KEYINPUT104), .A3(G868), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n831), .A2(new_n621), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(G295));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(G331));
  NAND2_X1  g482(.A1(new_n589), .A2(G168), .ZN(new_n908));
  NOR2_X1   g483(.A1(G171), .A2(G168), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n869), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G286), .B1(new_n586), .B2(new_n588), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n837), .B1(new_n912), .B2(new_n909), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n876), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n877), .A2(new_n882), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n911), .A2(new_n913), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n895), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n885), .ZN(new_n920));
  INV_X1    g495(.A(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(new_n922));
  INV_X1    g497(.A(new_n895), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n876), .B1(new_n919), .B2(new_n880), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n879), .A2(new_n881), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n911), .A2(new_n913), .A3(new_n927), .A4(KEYINPUT41), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n920), .B(new_n895), .C1(new_n921), .C2(new_n919), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  AND4_X1   g506(.A1(KEYINPUT43), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n918), .B2(new_n924), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n935), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT71), .B1(new_n471), .B2(new_n497), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n490), .A2(G126), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n509), .A2(new_n511), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n504), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G160), .A2(G40), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT107), .Z(new_n952));
  XNOR2_X1  g527(.A(new_n761), .B(new_n766), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n713), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1996), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n713), .A3(new_n957), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT106), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n808), .B(new_n811), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n814), .A2(new_n813), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT105), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n951), .C1(KEYINPUT105), .C2(new_n966), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n961), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n940), .C1(new_n943), .C2(new_n946), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n513), .B2(new_n940), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT50), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n975), .B(new_n474), .C1(new_n483), .C2(G2105), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n940), .C1(new_n943), .C2(new_n946), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n513), .A2(KEYINPUT115), .A3(new_n977), .A4(new_n940), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n974), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT120), .B(G1956), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n986));
  XNOR2_X1  g561(.A(G299), .B(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT110), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n513), .A2(new_n990), .A3(KEYINPUT45), .A4(new_n940), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n950), .B1(new_n948), .B2(new_n947), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(new_n444), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n985), .A2(new_n987), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n947), .A2(KEYINPUT111), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(new_n976), .A3(new_n971), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n998), .A2(new_n976), .A3(KEYINPUT122), .A4(new_n971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n766), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n977), .A3(new_n971), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n976), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1348), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n633), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n987), .B1(new_n985), .B2(new_n996), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n997), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT61), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n985), .A2(new_n987), .A3(new_n996), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(new_n1011), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT60), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1017));
  AOI21_X1  g592(.A(G2067), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1004), .A2(KEYINPUT60), .A3(new_n1009), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n619), .ZN(new_n1021));
  INV_X1    g596(.A(new_n987), .ZN(new_n1022));
  INV_X1    g597(.A(new_n984), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n998), .A2(new_n971), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n950), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(new_n982), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n989), .A2(new_n976), .A3(new_n949), .A4(new_n991), .ZN(new_n1027));
  INV_X1    g602(.A(new_n995), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1022), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n997), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1015), .A2(new_n1021), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT58), .B(G1341), .Z(new_n1033));
  NAND3_X1  g608(.A1(new_n1001), .A2(new_n1002), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT123), .B(G1996), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n992), .A2(new_n993), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n567), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT59), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1004), .A2(KEYINPUT60), .A3(new_n633), .A4(new_n1009), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n1040), .C1(new_n1037), .C2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1012), .B1(new_n1032), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT125), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT117), .B(G2084), .Z(new_n1045));
  NOR2_X1   g620(.A1(new_n950), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1005), .A2(new_n1006), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n948), .B1(new_n972), .B2(new_n973), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n976), .A2(new_n988), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1966), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G168), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n998), .B2(new_n971), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n976), .A2(new_n988), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n778), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(KEYINPUT125), .A3(new_n1047), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G168), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1054), .A2(KEYINPUT51), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(KEYINPUT126), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT126), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1053), .B1(new_n1057), .B2(new_n1047), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1054), .A2(KEYINPUT51), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1059), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2090), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n974), .A2(new_n982), .A3(new_n1076), .A4(new_n976), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1027), .A2(new_n795), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1053), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1072), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT116), .B(new_n1074), .C1(new_n1081), .C2(new_n1053), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n999), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G288), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT113), .B(G1976), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n599), .A2(new_n799), .A3(new_n600), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1092), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(G8), .A3(new_n999), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT52), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1090), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n950), .A2(G2090), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1005), .A2(new_n1100), .A3(new_n1101), .A4(new_n1006), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1078), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1005), .A2(new_n1006), .A3(new_n1101), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1053), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1099), .B1(new_n1106), .B2(new_n1075), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1083), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1007), .A2(new_n780), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1027), .B2(G2078), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(G2078), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1049), .A2(new_n1050), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n589), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n993), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n993), .A2(new_n1116), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n992), .A3(new_n1118), .A4(new_n1112), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1120), .B2(new_n589), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1120), .B2(G171), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1114), .A2(new_n589), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1121), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1043), .A2(new_n1071), .A3(new_n1108), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1059), .B(new_n1128), .C1(new_n1062), .C2(new_n1070), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1115), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1083), .A2(new_n1107), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1106), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1133), .A2(new_n1074), .A3(new_n1099), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1097), .A2(new_n1085), .A3(new_n788), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1084), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1126), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1133), .B2(new_n1074), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n1063), .B2(G286), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1067), .A2(new_n1143), .A3(G168), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1141), .A2(new_n1107), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1083), .A2(new_n1107), .A3(new_n1147), .A4(new_n1145), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n1140), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1083), .A2(new_n1107), .A3(new_n1145), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n969), .B1(new_n1139), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n951), .A2(new_n957), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n956), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n961), .A2(new_n964), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n951), .A2(new_n813), .A3(new_n814), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n808), .A2(new_n811), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n961), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(G2067), .B2(new_n761), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n952), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g741(.A1(G229), .A2(new_n463), .A3(G227), .ZN(new_n1168));
  NOR2_X1   g742(.A1(G401), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g743(.A(new_n1169), .B(new_n865), .C1(new_n936), .C2(new_n937), .ZN(G225));
  INV_X1    g744(.A(G225), .ZN(G308));
endmodule


