//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n467), .B1(new_n461), .B2(new_n462), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  AOI21_X1  g046(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n472));
  AOI22_X1  g047(.A1(G124), .A2(new_n472), .B1(new_n463), .B2(G136), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT70), .Z(G162));
  INV_X1    g054(.A(G138), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n481), .B(new_n486), .C1(new_n483), .C2(new_n482), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(KEYINPUT72), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT71), .A2(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT71), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(G126), .A2(new_n472), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n488), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n504), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  AOI22_X1  g087(.A1(new_n505), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n501), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  OR3_X1    g095(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n515), .B2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(G168));
  AOI22_X1  g098(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n503), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n506), .A2(new_n526), .B1(new_n508), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  AOI22_X1  g104(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n503), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n506), .A2(new_n533), .B1(new_n508), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT74), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(KEYINPUT76), .A3(new_n547), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n550), .B1(new_n545), .B2(KEYINPUT9), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n545), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n514), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n506), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(G651), .B1(new_n557), .B2(G91), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  OAI21_X1  g136(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n563));
  INV_X1    g138(.A(G87), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n506), .ZN(G288));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  INV_X1    g141(.A(G86), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n506), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n505), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G48), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n499), .B2(new_n500), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT78), .A4(G86), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n568), .A2(new_n570), .A3(new_n576), .A4(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n503), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n506), .A2(new_n581), .B1(new_n508), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT79), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n501), .A2(new_n505), .A3(G92), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n514), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n569), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT80), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G321));
  NOR2_X1   g172(.A1(G299), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g174(.A(new_n598), .B1(G868), .B2(G168), .ZN(G280));
  XNOR2_X1  g175(.A(KEYINPUT81), .B(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(G860), .B2(new_n601), .ZN(G148));
  NOR2_X1   g177(.A1(new_n536), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n601), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT82), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(G868), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n461), .A2(new_n462), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n465), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n463), .A2(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n472), .A2(G123), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n464), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n632), .B2(new_n634), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT17), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n642), .B2(new_n639), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  INV_X1    g223(.A(new_n639), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n645), .A3(new_n641), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n640), .A2(new_n645), .A3(new_n642), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  AOI211_X1 g240(.A(new_n663), .B(new_n665), .C1(new_n658), .C2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(G1981), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1971), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT33), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1976), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n684), .A2(KEYINPUT34), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT34), .B1(new_n684), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n674), .A2(G24), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n584), .B2(new_n674), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  OR2_X1    g268(.A1(G25), .A2(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n463), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n472), .A2(G119), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n464), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR4_X1   g279(.A1(new_n693), .A2(KEYINPUT89), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n689), .A2(new_n690), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  INV_X1    g285(.A(G28), .ZN(new_n711));
  AOI21_X1  g286(.A(G29), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n711), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT95), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n710), .B1(new_n713), .B2(new_n717), .C1(new_n619), .C2(new_n700), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(G29), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G160), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n674), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n537), .B2(new_n674), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n726), .B1(new_n725), .B2(new_n724), .C1(new_n728), .C2(G1341), .ZN(new_n729));
  NOR2_X1   g304(.A1(G27), .A2(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G164), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2078), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n674), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n674), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G1966), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n674), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n674), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n728), .A2(G1341), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n463), .A2(G139), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n608), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n464), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G2072), .Z(new_n748));
  NAND4_X1  g323(.A1(new_n733), .A2(new_n736), .A3(new_n740), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n674), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n595), .B2(new_n674), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n700), .A2(G35), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT98), .Z(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n700), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT29), .B(G2090), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n751), .A2(G1348), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n700), .A2(G32), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n472), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  OAI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(new_n700), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n752), .A2(new_n757), .A3(new_n758), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n739), .A2(new_n737), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n700), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n463), .A2(G140), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT90), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n472), .A2(G128), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n464), .A2(G116), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n771), .B(new_n783), .C1(G1966), .C2(new_n735), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n674), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n749), .A2(new_n769), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n708), .A2(new_n709), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(G311));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(G150));
  AOI22_X1  g369(.A1(new_n557), .A2(G93), .B1(new_n569), .B2(G55), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n503), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT100), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(new_n536), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n536), .A2(new_n797), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT38), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n595), .A2(G559), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n805));
  AOI21_X1  g380(.A(G860), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n798), .A2(G860), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT37), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(G145));
  XNOR2_X1  g385(.A(new_n610), .B(new_n699), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n472), .A2(G130), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT102), .ZN(new_n813));
  INV_X1    g388(.A(G118), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n814), .A2(KEYINPUT103), .A3(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT103), .B1(new_n814), .B2(G2105), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n815), .A2(new_n818), .B1(new_n463), .B2(G142), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n811), .B(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT104), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n781), .B(new_n497), .ZN(new_n823));
  INV_X1    g398(.A(new_n764), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n746), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n765), .B2(new_n746), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n823), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n822), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(G162), .B(new_n723), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n619), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  MUX2_X1   g408(.A(new_n821), .B(new_n822), .S(new_n827), .Z(new_n834));
  OAI211_X1 g409(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n831), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g411(.A(G868), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n798), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n605), .B(new_n801), .ZN(new_n839));
  INV_X1    g414(.A(new_n594), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G299), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(new_n841), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n839), .A2(KEYINPUT106), .A3(new_n846), .ZN(new_n850));
  INV_X1    g425(.A(new_n841), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n849), .B(new_n850), .C1(new_n839), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n584), .B(new_n680), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n854));
  XNOR2_X1  g429(.A(G303), .B(G305), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n852), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n838), .B1(new_n862), .B2(new_n837), .ZN(G295));
  OAI21_X1  g438(.A(new_n838), .B1(new_n862), .B2(new_n837), .ZN(G331));
  INV_X1    g439(.A(KEYINPUT109), .ZN(new_n865));
  XNOR2_X1  g440(.A(G168), .B(G301), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n801), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n799), .A2(new_n800), .A3(new_n866), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n841), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n859), .B(new_n870), .C1(new_n872), .C2(new_n845), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(new_n833), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n870), .B1(new_n872), .B2(new_n845), .ZN(new_n875));
  INV_X1    g450(.A(new_n859), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT43), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n871), .B1(new_n851), .B2(new_n842), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n841), .A2(KEYINPUT41), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n876), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n874), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n865), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g463(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n879), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n878), .A2(KEYINPUT43), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n874), .A2(new_n883), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT44), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n888), .A2(new_n889), .B1(new_n890), .B2(new_n892), .ZN(G397));
  INV_X1    g468(.A(KEYINPUT63), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n895));
  INV_X1    g470(.A(G1384), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n497), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n898));
  INV_X1    g473(.A(G2090), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT50), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n497), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n900), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n908));
  AOI21_X1  g483(.A(G1971), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n895), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n493), .A2(new_n495), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n472), .A2(G126), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n490), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G1384), .B1(new_n913), .B2(new_n488), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n901), .B1(new_n914), .B2(KEYINPUT45), .ZN(new_n915));
  INV_X1    g490(.A(new_n908), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(KEYINPUT110), .B(new_n904), .C1(new_n917), .C2(G1971), .ZN(new_n918));
  NAND2_X1  g493(.A1(G303), .A2(G8), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n910), .A2(new_n918), .A3(G8), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G8), .B1(new_n905), .B2(new_n909), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n901), .A2(new_n497), .A3(new_n896), .ZN(new_n925));
  INV_X1    g500(.A(G1976), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT52), .B1(G288), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n680), .A2(G1976), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n925), .A2(new_n927), .A3(G8), .A4(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT111), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT49), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n570), .A2(new_n576), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n506), .A2(new_n567), .ZN(new_n933));
  OAI21_X1  g508(.A(G1981), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(G305), .A2(G1981), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n914), .B2(new_n901), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n934), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n925), .A2(G8), .A3(new_n928), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT52), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n930), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n922), .A2(new_n924), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n497), .B2(new_n896), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n900), .ZN(new_n949));
  OAI211_X1 g524(.A(KEYINPUT112), .B(new_n901), .C1(new_n914), .C2(KEYINPUT45), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n908), .ZN(new_n951));
  INV_X1    g526(.A(G1966), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(KEYINPUT113), .A3(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n898), .A2(new_n901), .A3(new_n903), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n725), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT113), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  OAI211_X1 g532(.A(G8), .B(G168), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n894), .B1(new_n946), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n961), .B(new_n894), .C1(new_n946), .C2(new_n958), .ZN(new_n962));
  INV_X1    g537(.A(new_n958), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n910), .A2(new_n918), .A3(G8), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n894), .B1(new_n964), .B2(new_n920), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n922), .A3(new_n945), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n922), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n941), .A2(new_n926), .A3(new_n680), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G1981), .B2(G305), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n968), .A2(new_n945), .B1(new_n939), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n898), .A2(new_n901), .A3(new_n903), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n788), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(G2072), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n907), .A2(new_n908), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n553), .A2(new_n978), .A3(new_n558), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n553), .B2(new_n558), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1348), .ZN(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  INV_X1    g560(.A(new_n925), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n972), .A2(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n594), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n973), .A2(new_n976), .A3(new_n981), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n973), .A2(new_n981), .A3(new_n991), .A4(new_n976), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n986), .A2(new_n985), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT60), .B(new_n995), .C1(new_n954), .C2(G1348), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n594), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n954), .B2(G1348), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT60), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(KEYINPUT60), .A3(new_n840), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT58), .B(G1341), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n925), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n908), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1003), .B(new_n1005), .C1(new_n915), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n897), .A2(new_n906), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(new_n1006), .A3(new_n901), .A4(new_n908), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1003), .B1(new_n1011), .B2(new_n1005), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n537), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n537), .B(new_n1016), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n983), .A2(new_n989), .A3(KEYINPUT61), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1002), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT61), .B1(new_n993), .B2(new_n983), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n994), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  INV_X1    g598(.A(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1010), .A2(new_n1024), .A3(new_n901), .A4(new_n908), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1023), .A2(new_n1025), .B1(new_n972), .B2(new_n737), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n900), .B(KEYINPUT120), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(new_n948), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n900), .B(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n1010), .A3(KEYINPUT121), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1023), .A2(G2078), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1029), .A2(new_n1032), .A3(new_n908), .A4(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1026), .A2(G301), .A3(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n949), .A2(new_n950), .A3(new_n908), .A4(new_n1033), .ZN(new_n1036));
  AOI21_X1  g611(.A(G301), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1022), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT122), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1022), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT123), .B1(new_n1043), .B2(G171), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1026), .A2(G301), .A3(new_n1036), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT54), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n946), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1021), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n951), .A2(new_n952), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n955), .A3(new_n953), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G168), .A2(new_n938), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(KEYINPUT119), .B2(KEYINPUT51), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n1054), .B2(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n956), .B2(new_n957), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1057), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n967), .B(new_n971), .C1(new_n1050), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1056), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT62), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1056), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1037), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n946), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT125), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(new_n1080), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1072), .A2(new_n1021), .A3(new_n1042), .A4(new_n1049), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(KEYINPUT124), .A3(new_n967), .A4(new_n971), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1069), .A2(new_n1079), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1010), .A2(new_n900), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n781), .B(new_n985), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n765), .A2(new_n1006), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1086), .B(new_n1087), .C1(new_n1006), .C2(new_n824), .ZN(new_n1088));
  INV_X1    g663(.A(new_n702), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n699), .B(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n584), .B(G1986), .Z(new_n1093));
  OAI21_X1  g668(.A(new_n1085), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1085), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1086), .B2(new_n824), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT127), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1085), .A2(new_n1006), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT46), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT47), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n699), .B(new_n1089), .C1(new_n1088), .C2(new_n1085), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n781), .A2(G2067), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1103), .A2(KEYINPUT126), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT126), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1085), .A3(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1096), .A2(G1986), .A3(G290), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1108), .B(KEYINPUT48), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1096), .B2(new_n1091), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1095), .A2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g688(.A(new_n459), .ZN(new_n1115));
  NOR3_X1   g689(.A1(G229), .A2(new_n1115), .A3(G227), .ZN(new_n1116));
  INV_X1    g690(.A(G401), .ZN(new_n1117));
  NAND4_X1  g691(.A1(new_n1116), .A2(new_n835), .A3(new_n1117), .A4(new_n886), .ZN(G225));
  INV_X1    g692(.A(G225), .ZN(G308));
endmodule


