//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(KEYINPUT66), .A3(G101), .A4(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(G137), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n464), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n463), .A2(G136), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g057(.A(KEYINPUT68), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  INV_X1    g060(.A(G100), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n486), .A2(new_n464), .A3(KEYINPUT69), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n486), .B2(new_n464), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n479), .A2(new_n485), .A3(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n472), .B2(new_n473), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n464), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n472), .B2(new_n473), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n464), .C1(new_n460), .C2(new_n461), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT5), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n510), .B1(new_n506), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT71), .A3(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT70), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT70), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(KEYINPUT6), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n511), .A2(new_n517), .A3(G88), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(G543), .A3(new_n520), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n519), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n521), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n511), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n511), .A2(new_n517), .A3(G89), .A4(new_n520), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n517), .A2(G51), .A3(G543), .A4(new_n520), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G168));
  NAND4_X1  g111(.A1(new_n511), .A2(new_n517), .A3(G90), .A4(new_n520), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G52), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n517), .A2(G543), .A3(new_n520), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n506), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n508), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n541));
  NOR3_X1   g116(.A1(new_n506), .A2(KEYINPUT72), .A3(G543), .ZN(new_n542));
  OAI211_X1 g117(.A(G64), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n526), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n537), .B(new_n539), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR3_X1   g123(.A1(new_n548), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  NAND4_X1  g125(.A1(new_n517), .A2(G43), .A3(G543), .A4(new_n520), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n511), .A2(new_n517), .A3(G81), .A4(new_n520), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n526), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT76), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n511), .B2(G65), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n513), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n517), .A2(new_n520), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(G91), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n517), .A2(G53), .A3(G543), .A4(new_n520), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n569), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  NAND3_X1  g149(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G286));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n527), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n524), .A2(new_n526), .ZN(new_n578));
  INV_X1    g153(.A(new_n522), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G50), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT77), .A4(new_n521), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n577), .A2(new_n581), .ZN(G303));
  NAND4_X1  g157(.A1(new_n511), .A2(new_n517), .A3(G87), .A4(new_n520), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n517), .A2(G49), .A3(G543), .A4(new_n520), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n511), .A2(new_n517), .A3(G86), .A4(new_n520), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n522), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n511), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n526), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n587), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n592), .B1(new_n566), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n525), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n517), .A2(new_n520), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n598), .A2(G48), .A3(G543), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n597), .A2(new_n599), .A3(KEYINPUT78), .A4(new_n588), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n594), .A2(new_n600), .ZN(G305));
  NAND4_X1  g176(.A1(new_n517), .A2(G47), .A3(G543), .A4(new_n520), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n511), .A2(new_n517), .A3(G85), .A4(new_n520), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n526), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n511), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n513), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G54), .B2(new_n579), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n598), .A2(G91), .A3(new_n511), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n513), .B2(new_n563), .ZN(new_n621));
  INV_X1    g196(.A(new_n571), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n569), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n619), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n616), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n616), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT79), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g208(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n474), .A2(new_n464), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n643));
  OAI22_X1  g218(.A1(new_n640), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G123), .B2(new_n484), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n638), .A2(new_n639), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n651), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT17), .Z(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n665), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2096), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(G227));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  OR2_X1    g262(.A1(new_n680), .A2(new_n682), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n685), .A3(new_n683), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n689), .C1(new_n685), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT84), .B(G1986), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n700), .A3(new_n698), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n594), .A2(new_n600), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n706), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G6), .B2(new_n706), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT85), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G23), .B(G288), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n712), .A2(new_n714), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n705), .B1(new_n721), .B2(KEYINPUT34), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n705), .A3(KEYINPUT34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n484), .A2(G119), .ZN(new_n735));
  OR2_X1    g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n471), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n463), .A2(G131), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n730), .A2(new_n731), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n732), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n727), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n725), .A2(new_n726), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n706), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n555), .B2(new_n706), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n706), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G168), .B2(new_n706), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n750), .A2(G1341), .B1(G1966), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT91), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n733), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n761));
  INV_X1    g336(.A(G140), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n760), .A2(new_n761), .B1(new_n640), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G128), .B2(new_n484), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n733), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n753), .B(new_n766), .C1(G1341), .C2(new_n750), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n733), .B1(new_n768), .B2(G28), .ZN(new_n770));
  AND2_X1   g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NOR2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n645), .B2(G29), .ZN(new_n774));
  AND2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n733), .B1(KEYINPUT24), .B2(G34), .ZN(new_n776));
  OAI22_X1  g351(.A1(G160), .A2(new_n733), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT26), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(G141), .B(new_n464), .C1(new_n460), .C2(new_n461), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n484), .B2(G129), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(new_n733), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n733), .B2(G32), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n774), .B1(new_n777), .B2(G2084), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n733), .A2(G27), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT94), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n504), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n752), .A2(G1966), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n777), .A2(G2084), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n733), .A2(G33), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G139), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n640), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n464), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n799), .B1(new_n807), .B2(new_n733), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n798), .B1(G2072), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n797), .B(new_n809), .C1(G2072), .C2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n767), .A2(new_n796), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n733), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n733), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n814));
  INV_X1    g389(.A(G2090), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n813), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n612), .A2(new_n615), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G16), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n706), .A2(G4), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n817), .B1(G1348), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G5), .A2(G16), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT93), .Z(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G301), .B2(new_n706), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1961), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n788), .A2(new_n789), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT92), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n821), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n823), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n706), .A2(G20), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT23), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n624), .B2(new_n706), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1956), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n811), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n748), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n726), .B1(new_n725), .B2(new_n747), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(G311));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n748), .A3(new_n837), .ZN(G150));
  NOR2_X1   g417(.A1(new_n818), .A2(new_n627), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n517), .A2(G55), .A3(G543), .A4(new_n520), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n511), .A2(new_n517), .A3(G93), .A4(new_n520), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n526), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n555), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n554), .A2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n845), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT97), .B(G860), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n850), .A2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(G162), .B(G160), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n645), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n640), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G130), .B2(new_n484), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT100), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n635), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n740), .ZN(new_n872));
  INV_X1    g447(.A(new_n491), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n460), .B2(new_n461), .ZN(new_n874));
  AOI21_X1  g449(.A(G2105), .B1(new_n874), .B2(new_n493), .ZN(new_n875));
  OAI21_X1  g450(.A(G126), .B1(new_n460), .B2(new_n461), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n464), .B1(new_n876), .B2(new_n498), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G129), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n482), .B2(new_n483), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n878), .B(new_n503), .C1(new_n880), .C2(new_n785), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n484), .A2(G129), .ZN(new_n882));
  INV_X1    g457(.A(new_n785), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n504), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n881), .A2(new_n764), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n764), .B1(new_n881), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n807), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n484), .A2(G128), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n463), .A2(G140), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n890), .B(new_n891), .C1(new_n760), .C2(new_n761), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n504), .A2(new_n882), .A3(new_n883), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n786), .A2(new_n504), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(new_n884), .A3(new_n764), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(KEYINPUT98), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n807), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n887), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g475(.A(KEYINPUT99), .B(new_n807), .C1(new_n889), .C2(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n864), .B1(new_n872), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT101), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  INV_X1    g479(.A(new_n807), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT98), .B1(new_n895), .B2(new_n896), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT99), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n899), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n887), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n872), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT102), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n916), .B(new_n872), .C1(new_n904), .C2(new_n912), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n903), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n902), .B(new_n872), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n864), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  XNOR2_X1  g498(.A(new_n629), .B(new_n853), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n818), .A2(new_n624), .ZN(new_n925));
  NAND3_X1  g500(.A1(G299), .A2(new_n612), .A3(new_n615), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n925), .A2(KEYINPUT41), .A3(new_n926), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT41), .B1(new_n925), .B2(new_n926), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(new_n934), .A3(new_n927), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G288), .A2(KEYINPUT104), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n710), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n594), .A3(new_n600), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n527), .B(G290), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n947), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n937), .B2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(new_n938), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n929), .A2(new_n933), .A3(new_n953), .A4(new_n935), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n939), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n939), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n850), .A2(G868), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n958), .ZN(G331));
  OAI21_X1  g535(.A(G286), .B1(new_n547), .B2(new_n549), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n545), .A2(new_n546), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT73), .B1(new_n548), .B2(new_n526), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n537), .A2(new_n539), .ZN(new_n964));
  NAND4_X1  g539(.A1(G168), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n853), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n851), .A2(new_n961), .A3(new_n852), .A4(new_n965), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n930), .B2(new_n931), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(KEYINPUT106), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n853), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n554), .A2(new_n849), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n554), .A2(new_n849), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n961), .A4(new_n965), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n927), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n970), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n943), .A2(new_n947), .A3(new_n945), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n947), .B1(new_n943), .B2(new_n945), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n949), .A2(KEYINPUT108), .A3(new_n950), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G37), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n927), .A2(new_n967), .A3(new_n968), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n971), .A2(new_n973), .B1(new_n975), .B2(new_n980), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n951), .B(new_n993), .C1(new_n932), .C2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(new_n998), .A3(new_n992), .A4(new_n995), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n999), .A3(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n992), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n988), .A2(new_n989), .ZN(new_n1003));
  INV_X1    g578(.A(new_n931), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n982), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1003), .B1(new_n1007), .B2(new_n993), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n991), .A2(new_n1010), .A3(new_n992), .A4(new_n995), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1016), .B2(new_n1001), .ZN(new_n1017));
  AOI211_X1 g592(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(G397));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n469), .B(G40), .C1(new_n464), .C2(new_n475), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n504), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n878), .B2(new_n503), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1966), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1021), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1026), .A2(KEYINPUT113), .A3(new_n1031), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1032), .B(new_n1033), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1020), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT51), .B1(new_n1038), .B2(KEYINPUT124), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1037), .A3(G168), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(G286), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(G8), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1043), .B(KEYINPUT51), .C1(KEYINPUT124), .C2(new_n1038), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n577), .A2(new_n581), .A3(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1032), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1026), .A2(new_n1059), .A3(KEYINPUT45), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n1024), .B2(new_n1022), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1025), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1971), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1058), .A2(new_n815), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1054), .B(new_n1055), .C1(new_n1020), .C2(new_n1064), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1028), .A2(KEYINPUT125), .A3(G2078), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT125), .B1(new_n1028), .B2(G2078), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT53), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1062), .B2(G2078), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1032), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1071));
  INV_X1    g646(.A(G1961), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1051), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n1055), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1032), .B(new_n815), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1020), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n1020), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  OR2_X1    g660(.A1(G288), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1085), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n597), .A2(new_n599), .A3(new_n692), .A4(new_n588), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT49), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT115), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1094), .B(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1091), .B1(new_n1084), .B2(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1065), .A2(new_n1075), .A3(new_n1082), .A4(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1046), .A2(new_n1048), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G288), .A2(G1976), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT116), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1093), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1084), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1038), .A2(G168), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1065), .A2(new_n1098), .A3(new_n1082), .A4(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1038), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n1082), .A4(new_n1098), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1106), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n568), .B(new_n572), .C1(KEYINPUT118), .C2(KEYINPUT57), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n620), .B(KEYINPUT118), .C1(new_n513), .C2(new_n563), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1118), .B(new_n1119), .C1(new_n621), .C2(new_n623), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1025), .A2(new_n1060), .A3(new_n1061), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1116), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(KEYINPUT119), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1117), .A2(new_n1120), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT120), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1126), .A2(new_n1127), .A3(new_n1132), .A4(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G2067), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1071), .A2(new_n830), .B1(new_n1135), .B2(new_n1083), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(new_n818), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1125), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n818), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT121), .B(G1996), .Z(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT58), .B(G1341), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1062), .A2(new_n1142), .B1(new_n1083), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n554), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1136), .A2(new_n1139), .A3(new_n616), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1144), .B(new_n1145), .C1(KEYINPUT122), .C2(KEYINPUT59), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1126), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT61), .B1(new_n1152), .B2(new_n1124), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1141), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1125), .A2(KEYINPUT123), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1125), .A2(KEYINPUT123), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1134), .A2(new_n1155), .A3(KEYINPUT61), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1138), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1065), .A2(new_n1098), .A3(new_n1082), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n469), .A2(KEYINPUT53), .A3(G40), .A4(new_n794), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n475), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n464), .B1(new_n475), .B2(new_n1162), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1024), .A2(new_n1022), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1165), .A2(new_n1060), .A3(new_n1061), .A4(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1070), .A2(new_n1073), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(G171), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1160), .B1(new_n1075), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1068), .A2(new_n1074), .A3(G301), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1160), .B1(new_n1168), .B2(G171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1159), .A2(new_n1045), .A3(new_n1170), .A4(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1100), .B(new_n1114), .C1(new_n1158), .C2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1166), .A2(new_n1021), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n764), .B(G2067), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n786), .B(G1996), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n740), .B(new_n743), .Z(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n731), .B2(new_n728), .ZN(new_n1182));
  NOR2_X1   g757(.A1(G290), .A2(G1986), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT111), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1176), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1177), .B2(new_n786), .ZN(new_n1188));
  INV_X1    g763(.A(G1996), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1176), .A2(KEYINPUT46), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT46), .B1(new_n1176), .B2(new_n1189), .ZN(new_n1191));
  OR3_X1    g766(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT47), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n741), .A2(new_n743), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1179), .A2(new_n1195), .B1(G2067), .B2(new_n892), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1192), .A2(new_n1193), .B1(new_n1176), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT48), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1184), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1187), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1184), .A2(KEYINPUT48), .A3(new_n1176), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1200), .B(new_n1201), .C1(new_n1187), .C2(new_n1181), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1194), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1186), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g779(.A1(new_n918), .A2(new_n920), .ZN(new_n1206));
  OR3_X1    g780(.A1(G227), .A2(new_n458), .A3(G401), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n702), .B2(new_n703), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n1206), .A2(new_n1016), .A3(new_n1208), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


