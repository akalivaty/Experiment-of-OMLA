

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594;

  NOR2_X1 U328 ( .A1(n525), .A2(n468), .ZN(n469) );
  XNOR2_X1 U329 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n393) );
  XNOR2_X1 U330 ( .A(n317), .B(KEYINPUT84), .ZN(n318) );
  XOR2_X1 U331 ( .A(KEYINPUT13), .B(G57GAT), .Z(n367) );
  XNOR2_X1 U332 ( .A(n319), .B(n318), .ZN(n321) );
  OR2_X1 U333 ( .A1(n352), .A2(n351), .ZN(n353) );
  XNOR2_X1 U334 ( .A(n349), .B(n323), .ZN(n324) );
  XNOR2_X1 U335 ( .A(n394), .B(n393), .ZN(n418) );
  XNOR2_X1 U336 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U337 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U338 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U339 ( .A(n381), .B(n380), .Z(n587) );
  XNOR2_X1 U340 ( .A(n498), .B(n497), .ZN(n505) );
  XNOR2_X1 U341 ( .A(n452), .B(KEYINPUT58), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n297) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(KEYINPUT74), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U346 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n299) );
  XNOR2_X1 U347 ( .A(G190GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n312) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n302), .B(KEYINPUT8), .ZN(n343) );
  XOR2_X1 U352 ( .A(n343), .B(KEYINPUT64), .Z(n304) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U355 ( .A(G85GAT), .B(G92GAT), .Z(n351) );
  XOR2_X1 U356 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U357 ( .A(n351), .B(n423), .Z(n306) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G218GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U361 ( .A(G43GAT), .B(G134GAT), .Z(n439) );
  INV_X1 U362 ( .A(n439), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n562) );
  INV_X1 U365 ( .A(n562), .ZN(n478) );
  XNOR2_X1 U366 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n313), .B(KEYINPUT17), .ZN(n314) );
  XOR2_X1 U368 ( .A(n314), .B(KEYINPUT19), .Z(n316) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n447) );
  XNOR2_X1 U371 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n319) );
  INV_X1 U372 ( .A(KEYINPUT85), .ZN(n317) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n422) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G8GAT), .Z(n339) );
  XNOR2_X1 U376 ( .A(n422), .B(n339), .ZN(n325) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G204GAT), .Z(n322) );
  XNOR2_X1 U378 ( .A(G64GAT), .B(n322), .ZN(n349) );
  AND2_X1 U379 ( .A1(G226GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(G92GAT), .B(KEYINPUT90), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n447), .B(n328), .ZN(n464) );
  XOR2_X1 U383 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n429) );
  XNOR2_X1 U387 ( .A(G15GAT), .B(G1GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n331), .B(KEYINPUT71), .ZN(n368) );
  XOR2_X1 U389 ( .A(n429), .B(n368), .Z(n333) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n347) );
  XOR2_X1 U393 ( .A(KEYINPUT29), .B(G197GAT), .Z(n337) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G50GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U396 ( .A(n338), .B(G113GAT), .Z(n341) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(n339), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U399 ( .A(n342), .B(KEYINPUT72), .Z(n345) );
  XNOR2_X1 U400 ( .A(n343), .B(KEYINPUT67), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n507) );
  XNOR2_X1 U403 ( .A(G106GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n348), .B(G148GAT), .ZN(n424) );
  XNOR2_X1 U405 ( .A(n424), .B(n349), .ZN(n363) );
  XNOR2_X1 U406 ( .A(n367), .B(KEYINPUT31), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n350), .B(KEYINPUT73), .ZN(n352) );
  NAND2_X1 U408 ( .A1(n351), .A2(n352), .ZN(n354) );
  NAND2_X1 U409 ( .A1(n354), .A2(n353), .ZN(n356) );
  AND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n361) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G71GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n357), .B(G120GAT), .ZN(n442) );
  XNOR2_X1 U414 ( .A(n442), .B(KEYINPUT33), .ZN(n359) );
  INV_X1 U415 ( .A(KEYINPUT32), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n584) );
  XNOR2_X1 U417 ( .A(KEYINPUT41), .B(n584), .ZN(n508) );
  NOR2_X1 U418 ( .A1(n507), .A2(n508), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n364), .B(KEYINPUT46), .ZN(n382) );
  XOR2_X1 U420 ( .A(G155GAT), .B(G211GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G71GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n381) );
  XOR2_X1 U423 ( .A(n367), .B(G183GAT), .Z(n370) );
  XNOR2_X1 U424 ( .A(n368), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U426 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n372) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT14), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U431 ( .A(G8GAT), .B(G78GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n377), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U435 ( .A1(n382), .A2(n587), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n383), .B(KEYINPUT113), .ZN(n384) );
  NOR2_X1 U437 ( .A1(n384), .A2(n562), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n385), .B(KEYINPUT47), .ZN(n391) );
  XNOR2_X1 U439 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n387) );
  XNOR2_X1 U440 ( .A(KEYINPUT36), .B(n562), .ZN(n590) );
  NAND2_X1 U441 ( .A1(n587), .A2(n590), .ZN(n386) );
  XOR2_X1 U442 ( .A(n387), .B(n386), .Z(n388) );
  NOR2_X1 U443 ( .A1(n584), .A2(n388), .ZN(n389) );
  NAND2_X1 U444 ( .A1(n389), .A2(n507), .ZN(n390) );
  NAND2_X1 U445 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n392), .B(KEYINPUT48), .ZN(n554) );
  NAND2_X1 U447 ( .A1(n464), .A2(n554), .ZN(n394) );
  XOR2_X1 U448 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n396) );
  XNOR2_X1 U449 ( .A(G141GAT), .B(G148GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n405) );
  XOR2_X1 U451 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n403) );
  XOR2_X1 U452 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n398) );
  XNOR2_X1 U453 ( .A(KEYINPUT77), .B(G127GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(G113GAT), .B(n399), .Z(n448) );
  XOR2_X1 U456 ( .A(G155GAT), .B(KEYINPUT2), .Z(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n425) );
  XNOR2_X1 U459 ( .A(n448), .B(n425), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n417) );
  NAND2_X1 U462 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XOR2_X1 U463 ( .A(G162GAT), .B(G134GAT), .Z(n407) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G120GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT74), .B(G85GAT), .Z(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U469 ( .A(G57GAT), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n525) );
  NOR2_X1 U474 ( .A1(n418), .A2(n525), .ZN(n576) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n420) );
  XNOR2_X1 U476 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n433) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n431) );
  XOR2_X1 U480 ( .A(n425), .B(KEYINPUT24), .Z(n427) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n472) );
  NAND2_X1 U486 ( .A1(n576), .A2(n472), .ZN(n435) );
  XNOR2_X1 U487 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n451) );
  XOR2_X1 U489 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n437) );
  XNOR2_X1 U490 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT81), .Z(n441) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U495 ( .A(n442), .B(KEYINPUT79), .Z(n444) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n538) );
  NAND2_X1 U501 ( .A1(n451), .A2(n538), .ZN(n572) );
  NOR2_X1 U502 ( .A1(n478), .A2(n572), .ZN(n454) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n452) );
  NOR2_X1 U504 ( .A1(n507), .A2(n572), .ZN(n457) );
  INV_X1 U505 ( .A(G169GAT), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT120), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(n456), .ZN(G1348GAT) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U509 ( .A1(n538), .A2(n464), .ZN(n458) );
  XOR2_X1 U510 ( .A(KEYINPUT95), .B(n458), .Z(n459) );
  NAND2_X1 U511 ( .A1(n472), .A2(n459), .ZN(n461) );
  INV_X1 U512 ( .A(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(n466) );
  XNOR2_X1 U514 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n538), .A2(n472), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n463), .B(n462), .ZN(n577) );
  XNOR2_X1 U517 ( .A(KEYINPUT27), .B(n464), .ZN(n470) );
  NAND2_X1 U518 ( .A1(n577), .A2(n470), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U520 ( .A(KEYINPUT96), .B(n467), .Z(n468) );
  XNOR2_X1 U521 ( .A(KEYINPUT97), .B(n469), .ZN(n477) );
  XOR2_X1 U522 ( .A(n538), .B(KEYINPUT83), .Z(n474) );
  NAND2_X1 U523 ( .A1(n470), .A2(n525), .ZN(n471) );
  XNOR2_X1 U524 ( .A(n471), .B(KEYINPUT91), .ZN(n552) );
  XNOR2_X1 U525 ( .A(n472), .B(KEYINPUT28), .ZN(n490) );
  NAND2_X1 U526 ( .A1(n552), .A2(n490), .ZN(n539) );
  XNOR2_X1 U527 ( .A(n539), .B(KEYINPUT92), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U529 ( .A(KEYINPUT93), .B(n475), .ZN(n476) );
  NAND2_X1 U530 ( .A1(n477), .A2(n476), .ZN(n493) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n480) );
  NAND2_X1 U532 ( .A1(n587), .A2(n478), .ZN(n479) );
  XNOR2_X1 U533 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U534 ( .A1(n493), .A2(n481), .ZN(n482) );
  XNOR2_X1 U535 ( .A(n482), .B(KEYINPUT98), .ZN(n510) );
  NOR2_X1 U536 ( .A1(n507), .A2(n584), .ZN(n496) );
  INV_X1 U537 ( .A(n496), .ZN(n483) );
  NOR2_X1 U538 ( .A1(n510), .A2(n483), .ZN(n491) );
  NAND2_X1 U539 ( .A1(n525), .A2(n491), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n464), .A2(n491), .ZN(n486) );
  XNOR2_X1 U542 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U544 ( .A1(n491), .A2(n538), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  INV_X1 U547 ( .A(n490), .ZN(n533) );
  NAND2_X1 U548 ( .A1(n491), .A2(n533), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U551 ( .A1(n590), .A2(n493), .ZN(n494) );
  NOR2_X1 U552 ( .A1(n587), .A2(n494), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n495), .Z(n522) );
  NAND2_X1 U554 ( .A1(n522), .A2(n496), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT100), .B(KEYINPUT38), .Z(n497) );
  NAND2_X1 U556 ( .A1(n505), .A2(n525), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n505), .A2(n464), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n503) );
  NAND2_X1 U561 ( .A1(n505), .A2(n538), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n505), .A2(n533), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n512) );
  INV_X1 U567 ( .A(n507), .ZN(n579) );
  XNOR2_X1 U568 ( .A(n508), .B(KEYINPUT102), .ZN(n566) );
  NOR2_X1 U569 ( .A1(n579), .A2(n566), .ZN(n523) );
  INV_X1 U570 ( .A(n523), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n510), .A2(n509), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n525), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n464), .A2(n517), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(KEYINPUT104), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n538), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n533), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT105), .Z(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n524), .B(KEYINPUT107), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n534), .A2(n525), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT108), .ZN(n527) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  XOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT109), .Z(n529) );
  NAND2_X1 U591 ( .A1(n534), .A2(n464), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n534), .A2(n538), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT111), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n554), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(KEYINPUT114), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n549), .A2(n579), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U606 ( .A(n549), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n543), .A2(n566), .ZN(n545) );
  XNOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NAND2_X1 U611 ( .A1(n549), .A2(n587), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n562), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n556) );
  AND2_X1 U618 ( .A1(n577), .A2(n552), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n557) );
  INV_X1 U620 ( .A(n557), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n563), .A2(n579), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  NOR2_X1 U623 ( .A1(n508), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n587), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT117), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n572), .A2(n566), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  INV_X1 U638 ( .A(n587), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n578), .B(KEYINPUT124), .Z(n589) );
  AND2_X1 U644 ( .A1(n589), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n589), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n589), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n594) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(G1355GAT) );
endmodule

