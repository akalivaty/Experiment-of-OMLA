//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT74), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G15gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G113gat), .B2(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n217));
  OAI21_X1  g016(.A(G113gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n213), .A2(KEYINPUT71), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n210), .A2(new_n211), .B1(new_n213), .B2(KEYINPUT71), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n218), .A2(new_n208), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT25), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G183gat), .B(G190gat), .Z(new_n232));
  NOR3_X1   g031(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n232), .A2(KEYINPUT24), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n236), .A3(new_n225), .A4(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n229), .A2(new_n230), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n239), .B(new_n224), .C1(new_n225), .C2(KEYINPUT25), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n235), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n241), .A2(new_n223), .B1(new_n242), .B2(new_n233), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT27), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G183gat), .ZN(new_n249));
  INV_X1    g048(.A(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT28), .B1(new_n251), .B2(KEYINPUT66), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n250), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(KEYINPUT28), .A3(new_n250), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n252), .A2(new_n256), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n261), .A2(new_n266), .A3(new_n262), .A4(new_n263), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n239), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n222), .B(new_n245), .C1(new_n260), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n271), .B(new_n273), .C1(new_n257), .C2(new_n259), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n278), .A2(KEYINPUT72), .A3(new_n222), .A4(new_n245), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n245), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n215), .A2(new_n221), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n207), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n283), .B2(new_n285), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  AOI221_X4 g092(.A(new_n290), .B1(new_n287), .B2(new_n206), .C1(new_n283), .C2(new_n285), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n222), .B1(new_n278), .B2(new_n245), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n276), .B2(new_n275), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n284), .A4(new_n279), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n277), .A2(new_n282), .A3(new_n284), .A4(new_n279), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT77), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT34), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n284), .B2(KEYINPUT76), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n302), .ZN(new_n306));
  INV_X1    g105(.A(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n296), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n305), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n304), .B1(new_n300), .B2(new_n302), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n293), .B(new_n295), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT78), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n287), .B1(new_n283), .B2(new_n285), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n291), .A2(new_n315), .A3(new_n207), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(new_n294), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(new_n305), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n309), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT92), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(KEYINPUT78), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n314), .A3(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n309), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n280), .A2(KEYINPUT79), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n278), .A2(new_n328), .A3(new_n245), .ZN(new_n329));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336));
  INV_X1    g135(.A(G211gat), .ZN(new_n337));
  INV_X1    g136(.A(G218gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n340), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n278), .A2(new_n331), .A3(new_n245), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n333), .A2(new_n334), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n333), .A2(new_n344), .A3(new_n345), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT80), .ZN(new_n348));
  INV_X1    g147(.A(new_n329), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n328), .B1(new_n278), .B2(new_n245), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n331), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n280), .A2(new_n332), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n346), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n327), .A2(new_n329), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n331), .B1(new_n280), .B2(new_n332), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT80), .B(new_n347), .C1(new_n360), .C2(new_n344), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n346), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(KEYINPUT30), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n354), .A2(new_n365), .A3(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(G155gat), .B2(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(KEYINPUT82), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G141gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n388), .A3(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n379), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n383), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n376), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n343), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n384), .A2(new_n377), .B1(new_n390), .B2(new_n392), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n340), .A2(new_n342), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n341), .B1(new_n339), .B2(new_n335), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT87), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT87), .B(new_n406), .C1(new_n397), .C2(new_n402), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(G22gat), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(G228gat), .A3(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n407), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n371), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n410), .B2(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n412), .B(new_n371), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT89), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n412), .A2(new_n371), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n415), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n413), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(G57gat), .B(G85gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT83), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n385), .A2(new_n393), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n281), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n385), .A2(new_n393), .B1(new_n215), .B2(new_n221), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n222), .B1(KEYINPUT3), .B2(new_n433), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n432), .B1(new_n438), .B2(new_n395), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n222), .A2(new_n398), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n222), .A2(new_n398), .A3(KEYINPUT84), .A4(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT4), .B1(new_n433), .B2(new_n281), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n437), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n441), .A3(KEYINPUT85), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n449), .A3(new_n440), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n433), .A2(KEYINPUT3), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(new_n395), .A3(new_n281), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n454));
  INV_X1    g253(.A(new_n432), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n430), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n459));
  NAND4_X1  g258(.A1(new_n439), .A2(new_n454), .A3(new_n450), .A4(new_n448), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n453), .A2(new_n455), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n444), .A2(new_n445), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n443), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n460), .B(new_n429), .C1(new_n463), .C2(new_n437), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT91), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n458), .A2(new_n459), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n458), .A2(new_n464), .A3(new_n468), .A4(new_n459), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n367), .A2(new_n425), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n321), .A2(new_n326), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n465), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n364), .B2(new_n366), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n318), .B1(new_n296), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n424), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n324), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n448), .A2(new_n453), .A3(new_n450), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n432), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(KEYINPUT39), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n434), .A2(new_n435), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(KEYINPUT39), .C1(new_n432), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n488), .A3(new_n429), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT40), .A4(new_n429), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(new_n458), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n364), .A2(new_n366), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT90), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n362), .B1(new_n361), .B2(new_n346), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n470), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n360), .A2(new_n343), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n333), .A2(new_n345), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n343), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n354), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n502), .B(new_n362), .C1(new_n503), .C2(KEYINPUT37), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n362), .A2(KEYINPUT37), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n503), .A2(KEYINPUT37), .B1(new_n363), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n497), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n364), .A2(new_n493), .A3(new_n509), .A4(new_n366), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n508), .A3(new_n480), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n475), .A2(new_n480), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n324), .A2(new_n479), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n324), .A2(new_n516), .A3(new_n309), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n511), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n483), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G127gat), .B(G155gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT100), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n534), .B(new_n538), .C1(new_n535), .C2(G1gat), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(G15gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(G22gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n411), .A2(G15gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n536), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G8gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n537), .A2(new_n546), .B1(new_n548), .B2(KEYINPUT97), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(KEYINPUT97), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n549), .B(new_n550), .C1(new_n525), .C2(new_n524), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n531), .A2(new_n532), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n531), .A2(new_n532), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n550), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561));
  NAND2_X1  g360(.A1(G43gat), .A2(G50gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT95), .B(G43gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(G50gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  AND2_X1   g364(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G50gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n205), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n561), .B1(new_n574), .B2(new_n562), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n575), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT17), .B1(new_n576), .B2(new_n578), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT96), .B(KEYINPUT17), .Z(new_n583));
  OAI211_X1 g382(.A(new_n577), .B(new_n583), .C1(new_n572), .C2(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n580), .B(new_n581), .C1(new_n585), .C2(new_n560), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT99), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT18), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT18), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(KEYINPUT99), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n560), .B(new_n579), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n581), .B(KEYINPUT13), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G113gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n380), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT12), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n590), .A3(new_n593), .A4(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT7), .ZN(new_n610));
  INV_X1    g409(.A(G99gat), .ZN(new_n611));
  INV_X1    g410(.A(G106gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT8), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT101), .B(G85gat), .Z(new_n614));
  OAI211_X1 g413(.A(new_n610), .B(new_n613), .C1(G92gat), .C2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n524), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(new_n616), .ZN(new_n620));
  INV_X1    g419(.A(new_n524), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT10), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n608), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n622), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(new_n608), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  OR2_X1    g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n624), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n607), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n608), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n579), .A2(new_n620), .B1(KEYINPUT41), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n582), .A2(new_n584), .A3(new_n617), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n638), .A2(new_n639), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n640), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR4_X1   g451(.A1(new_n559), .A2(new_n606), .A3(new_n636), .A4(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n519), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n474), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(G1gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1324gat));
  INV_X1    g456(.A(new_n654), .ZN(new_n658));
  OAI21_X1  g457(.A(G8gat), .B1(new_n658), .B2(new_n367), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(new_n367), .ZN(new_n661));
  NAND2_X1  g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n535), .A2(new_n540), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n654), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n664), .A2(KEYINPUT104), .A3(new_n660), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT104), .B1(new_n664), .B2(new_n660), .ZN(new_n666));
  OAI221_X1 g465(.A(new_n659), .B1(new_n660), .B2(new_n664), .C1(new_n665), .C2(new_n666), .ZN(G1325gat));
  AND3_X1   g466(.A1(new_n324), .A2(new_n516), .A3(new_n309), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n516), .B1(new_n324), .B2(new_n479), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n658), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n321), .A2(new_n326), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n654), .A2(new_n542), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n424), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(new_n652), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n483), .B2(new_n518), .ZN(new_n680));
  INV_X1    g479(.A(new_n559), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(new_n606), .A3(new_n636), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n569), .A3(new_n474), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n682), .B(KEYINPUT105), .Z(new_n686));
  XOR2_X1   g485(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n519), .A2(new_n652), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n680), .A2(KEYINPUT108), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n680), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n668), .A2(new_n669), .A3(new_n512), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n696), .A2(new_n511), .B1(new_n472), .B2(new_n482), .ZN(new_n697));
  OAI211_X1 g496(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n697), .C2(new_n679), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n686), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(new_n474), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n685), .B1(new_n701), .B2(new_n569), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n565), .A3(new_n661), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  AND2_X1   g503(.A1(new_n700), .A2(new_n661), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n565), .ZN(G1329gat));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  INV_X1    g506(.A(new_n563), .ZN(new_n708));
  INV_X1    g507(.A(new_n670), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n683), .A2(new_n673), .A3(new_n708), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n711), .B(KEYINPUT109), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n670), .B(new_n686), .C1(new_n692), .C2(new_n699), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n715), .B(KEYINPUT47), .C1(new_n716), .C2(new_n708), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(G1330gat));
  NOR2_X1   g517(.A1(new_n480), .A2(G50gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n683), .A2(new_n719), .ZN(new_n720));
  AOI211_X1 g519(.A(new_n480), .B(new_n686), .C1(new_n692), .C2(new_n699), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT48), .B(new_n720), .C1(new_n721), .C2(new_n573), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(KEYINPUT110), .A3(new_n719), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n700), .A2(new_n424), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(G50gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n728), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g528(.A1(new_n681), .A2(new_n606), .A3(new_n679), .ZN(new_n730));
  INV_X1    g529(.A(new_n636), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT111), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n519), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n473), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g535(.A(new_n734), .B(KEYINPUT112), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n661), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT49), .B(G64gat), .Z(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n737), .A2(G71gat), .A3(new_n709), .ZN(new_n742));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n734), .B2(new_n672), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n424), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT113), .B(G78gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1335gat));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n519), .A2(new_n652), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n681), .A2(new_n605), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n680), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n731), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n614), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n474), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n636), .ZN(new_n759));
  AOI211_X1 g558(.A(new_n473), .B(new_n759), .C1(new_n692), .C2(new_n699), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n614), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n692), .B2(new_n699), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n763), .A2(new_n761), .A3(new_n474), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n762), .B2(new_n764), .ZN(G1336gat));
  INV_X1    g564(.A(G92gat), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n661), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n367), .A2(G92gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n367), .B(new_n759), .C1(new_n692), .C2(new_n699), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n769), .B(new_n772), .C1(new_n773), .C2(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1337gat));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n611), .A3(new_n673), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n763), .A2(new_n709), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n611), .ZN(G1338gat));
  AOI21_X1  g577(.A(new_n612), .B1(new_n763), .B2(new_n424), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n480), .A2(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT53), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n480), .B(new_n759), .C1(new_n692), .C2(new_n699), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n781), .B(new_n784), .C1(new_n785), .C2(new_n612), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n623), .A2(new_n624), .A3(new_n608), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n630), .B1(new_n625), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n635), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT55), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n790), .A2(new_n792), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(KEYINPUT115), .A3(new_n635), .A4(new_n793), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n800), .A3(new_n605), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n585), .A2(new_n560), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n581), .B1(new_n802), .B2(new_n580), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n591), .A2(new_n592), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n600), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n604), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n636), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n652), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n806), .A2(new_n652), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n809), .A2(new_n796), .A3(new_n800), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n559), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n730), .A2(new_n636), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n480), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n672), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n661), .A2(new_n473), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(KEYINPUT116), .A3(new_n480), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n210), .A3(new_n606), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n424), .B(new_n514), .C1(new_n811), .C2(new_n813), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n818), .ZN(new_n823));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n605), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(new_n824), .ZN(G1340gat));
  OAI21_X1  g624(.A(G120gat), .B1(new_n820), .B2(new_n731), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n216), .A2(new_n217), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(new_n827), .A3(new_n636), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1341gat));
  OAI21_X1  g628(.A(G127gat), .B1(new_n820), .B2(new_n559), .ZN(new_n830));
  INV_X1    g629(.A(G127gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n823), .A2(new_n831), .A3(new_n681), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1342gat));
  NOR2_X1   g632(.A1(new_n679), .A2(G134gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n822), .A2(new_n818), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT56), .Z(new_n836));
  NAND4_X1  g635(.A1(new_n817), .A2(new_n652), .A3(new_n818), .A4(new_n819), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n837), .B2(G134gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT118), .B(new_n836), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n670), .A2(new_n818), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n794), .A2(new_n795), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n807), .A2(new_n848), .B1(new_n849), .B2(new_n605), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n848), .B2(new_n807), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n810), .B1(new_n851), .B2(new_n679), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n813), .B1(new_n852), .B2(new_n681), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n480), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n480), .B1(new_n811), .B2(new_n813), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(KEYINPUT57), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n854), .B1(new_n853), .B2(new_n856), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n386), .ZN(new_n862));
  INV_X1    g661(.A(new_n388), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n861), .A2(new_n606), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n858), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n380), .A3(new_n605), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(G148gat), .C1(new_n861), .C2(new_n731), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n679), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n809), .A2(new_n849), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n681), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n855), .B(new_n424), .C1(new_n877), .C2(new_n812), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(new_n636), .C1(new_n855), .C2(new_n858), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n378), .B1(new_n880), .B2(new_n847), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n378), .A3(new_n636), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n861), .B2(new_n559), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n865), .A2(G155gat), .A3(new_n559), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n861), .A2(new_n892), .A3(new_n679), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n865), .B2(new_n679), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n815), .A2(new_n816), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n367), .A2(new_n474), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n673), .A3(new_n819), .A4(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n817), .A2(KEYINPUT122), .A3(new_n819), .A4(new_n897), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(G169gat), .A3(new_n605), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n822), .A2(new_n897), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n262), .B1(new_n903), .B2(new_n606), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n902), .A2(new_n904), .ZN(G1348gat));
  INV_X1    g704(.A(new_n903), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n263), .A3(new_n636), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n900), .A2(new_n636), .A3(new_n901), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n263), .ZN(G1349gat));
  NAND2_X1  g708(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n681), .A2(new_n254), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n681), .A3(new_n901), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(G183gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n915), .B(new_n912), .C1(new_n913), .C2(G183gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n250), .A3(new_n652), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n652), .A3(new_n901), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(G190gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n921), .B2(G190gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n814), .A2(new_n473), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n670), .A2(new_n661), .A3(new_n424), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(new_n927), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n605), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n878), .B1(new_n855), .B2(new_n858), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n670), .A2(new_n897), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n605), .A2(G197gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n731), .A2(G204gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n929), .A2(new_n930), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n929), .A2(KEYINPUT125), .A3(new_n930), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n939), .B1(new_n945), .B2(KEYINPUT62), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n943), .A2(KEYINPUT126), .A3(new_n947), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n879), .A2(new_n935), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n945), .A2(KEYINPUT62), .B1(new_n950), .B2(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n337), .A3(new_n681), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n681), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n932), .A2(new_n338), .A3(new_n652), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n934), .A2(new_n679), .A3(new_n935), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n338), .ZN(G1355gat));
endmodule


