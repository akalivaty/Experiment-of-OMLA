//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT71), .B(G218gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT72), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT22), .B1(new_n205), .B2(G211gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(new_n204), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n203), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n202), .B1(new_n208), .B2(KEYINPUT72), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G183gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G190gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n216), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n219), .A3(KEYINPUT28), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(KEYINPUT26), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(KEYINPUT26), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G169gat), .ZN(new_n235));
  INV_X1    g034(.A(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  OAI22_X1  g038(.A1(new_n235), .A2(new_n237), .B1(new_n239), .B2(new_n227), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n234), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n230), .A2(KEYINPUT23), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n238), .A2(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n228), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n244), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  INV_X1    g051(.A(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n255));
  AOI21_X1  g054(.A(G183gat), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n250), .B(KEYINPUT25), .C1(new_n251), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G169gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n248), .B1(new_n228), .B2(new_n247), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n242), .B(new_n244), .C1(G183gat), .C2(G190gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT25), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n256), .A2(new_n251), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n236), .A3(KEYINPUT23), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT25), .B(new_n269), .C1(new_n239), .C2(new_n227), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT66), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n246), .A2(new_n273), .A3(new_n257), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n223), .A2(new_n224), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n272), .A2(new_n274), .B1(new_n275), .B2(new_n232), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n215), .B(new_n260), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n246), .A2(new_n273), .A3(new_n257), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n246), .B2(new_n257), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n233), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n215), .A4(new_n260), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n215), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n233), .B(new_n259), .C1(new_n281), .C2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n278), .B1(new_n233), .B2(new_n258), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G8gat), .B(G36gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n287), .A2(KEYINPUT76), .A3(new_n292), .A4(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n280), .A2(new_n292), .A3(new_n286), .A4(new_n297), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n215), .B1(new_n290), .B2(new_n291), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n288), .A3(new_n260), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT37), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT84), .B(KEYINPUT37), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n280), .A2(new_n292), .A3(new_n286), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n297), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT38), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n302), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n287), .A2(new_n292), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n312), .A2(KEYINPUT37), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT38), .B1(new_n313), .B2(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT77), .ZN(new_n317));
  INV_X1    g116(.A(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT78), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT78), .B1(new_n319), .B2(new_n321), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n315), .B(new_n317), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n319), .A2(new_n321), .ZN(new_n327));
  INV_X1    g126(.A(new_n315), .ZN(new_n328));
  NOR3_X1   g127(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n332));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT68), .B1(new_n336), .B2(G113gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G113gat), .B2(new_n336), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n334), .B(new_n335), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(KEYINPUT1), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n344), .A3(new_n330), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n332), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n331), .B2(new_n343), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n326), .A2(new_n330), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n340), .A2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT4), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g153(.A(new_n347), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n331), .A2(new_n343), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n330), .A2(new_n326), .B1(new_n340), .B2(new_n342), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n359), .A3(KEYINPUT79), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(G85gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n362), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n353), .A2(new_n359), .A3(KEYINPUT79), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n359), .B1(KEYINPUT79), .B2(new_n353), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n366), .B(KEYINPUT83), .Z(new_n373));
  NAND3_X1  g172(.A1(new_n361), .A2(new_n362), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n311), .A2(new_n314), .A3(new_n367), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n298), .A2(new_n377), .A3(new_n301), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n312), .A2(new_n308), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n299), .A2(new_n377), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n356), .A2(new_n355), .A3(new_n357), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n346), .A2(new_n349), .A3(new_n352), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n355), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT39), .ZN(new_n385));
  INV_X1    g184(.A(new_n373), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n355), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n385), .B(new_n386), .C1(KEYINPUT39), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n381), .A2(new_n374), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT31), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G50gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n213), .B2(new_n214), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n344), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n331), .ZN(new_n399));
  INV_X1    g198(.A(G228gat), .ZN(new_n400));
  INV_X1    g199(.A(G233gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n345), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n215), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n399), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n350), .B1(new_n397), .B2(new_n344), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n215), .A2(new_n406), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n403), .B(new_n402), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n411), .A3(G22gat), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n408), .A2(new_n411), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT82), .B(G22gat), .Z(new_n414));
  OAI211_X1 g213(.A(new_n395), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n395), .B(KEYINPUT80), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n408), .A2(new_n414), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n408), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n376), .A2(new_n392), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n283), .A2(new_n351), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n233), .B(new_n343), .C1(new_n281), .C2(new_n282), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n426), .A3(new_n424), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  INV_X1    g233(.A(G71gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G99gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n438), .A3(new_n430), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n432), .A2(new_n433), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(KEYINPUT33), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n440), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n440), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n428), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n437), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n438), .B1(new_n429), .B2(new_n430), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n449), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n445), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n441), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n440), .A2(new_n442), .A3(new_n445), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n427), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n361), .A2(new_n362), .A3(new_n366), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n371), .A2(new_n372), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n367), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n420), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n455), .A3(KEYINPUT36), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n422), .A2(new_n458), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n420), .B1(new_n448), .B2(new_n455), .ZN(new_n467));
  INV_X1    g266(.A(new_n462), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n375), .A2(new_n367), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n456), .A2(new_n472), .A3(new_n421), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n465), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G29gat), .ZN(new_n475));
  INV_X1    g274(.A(G36gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT14), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(G29gat), .B2(G36gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT86), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n486), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT15), .B(new_n487), .C1(KEYINPUT87), .C2(new_n483), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n482), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n481), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(KEYINPUT17), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(G1gat), .ZN(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT16), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(KEYINPUT88), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n501), .A3(G8gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n492), .A2(KEYINPUT17), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n489), .A2(new_n491), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n507), .B2(new_n512), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n510), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n511), .A4(new_n510), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n515), .A2(new_n516), .B1(new_n512), .B2(new_n507), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n511), .B(KEYINPUT13), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT11), .B(G169gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XOR2_X1   g327(.A(G113gat), .B(G141gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT85), .Z(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT12), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n519), .A2(new_n534), .A3(new_n522), .A4(new_n525), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n474), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT92), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT41), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n541), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT95), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n493), .A2(new_n509), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n554), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n540), .ZN(new_n561));
  XOR2_X1   g360(.A(G134gat), .B(G162gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n558), .A2(new_n565), .A3(new_n559), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n560), .A2(KEYINPUT96), .A3(new_n563), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G64gat), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n571), .A2(G57gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(G57gat), .ZN(new_n573));
  AND2_X1   g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n572), .A2(new_n573), .B1(KEYINPUT9), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n507), .B1(KEYINPUT21), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT91), .Z(new_n579));
  XOR2_X1   g378(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n582));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n581), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n554), .A2(KEYINPUT10), .A3(new_n577), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n552), .B(new_n577), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G230gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n401), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n592), .A2(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n236), .ZN(new_n603));
  INV_X1    g402(.A(G204gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n599), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n598), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n612), .B2(new_n605), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n590), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n537), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n461), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT98), .B(G1gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(G1324gat));
  INV_X1    g418(.A(new_n381), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT42), .Z(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n503), .B2(new_n621), .ZN(G1325gat));
  INV_X1    g424(.A(new_n616), .ZN(new_n626));
  AOI21_X1  g425(.A(G15gat), .B1(new_n626), .B2(new_n456), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n458), .A2(new_n464), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(G15gat), .B2(new_n630), .ZN(G1326gat));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n421), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT43), .B(G22gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1327gat));
  NOR3_X1   g433(.A1(new_n568), .A2(new_n564), .A3(new_n566), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n474), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n589), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n613), .ZN(new_n638));
  INV_X1    g437(.A(new_n536), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n461), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n475), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT45), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n635), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n469), .B2(new_n473), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n467), .A2(new_n472), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n420), .B(new_n462), .C1(new_n455), .C2(new_n448), .ZN(new_n651));
  OAI211_X1 g450(.A(KEYINPUT100), .B(new_n650), .C1(new_n651), .C2(new_n466), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n465), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n649), .A2(new_n652), .A3(KEYINPUT101), .A4(new_n465), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n646), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n536), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n533), .A2(KEYINPUT99), .A3(new_n535), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n659), .A2(new_n638), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n643), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n645), .B1(new_n667), .B2(new_n475), .ZN(G1328gat));
  AOI21_X1  g467(.A(G36gat), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n642), .A2(new_n381), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n381), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n674), .B2(new_n476), .ZN(G1329gat));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  INV_X1    g475(.A(new_n456), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n486), .B1(new_n641), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n638), .A2(new_n664), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n628), .B(new_n679), .C1(new_n657), .C2(new_n658), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(new_n486), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n685), .B(new_n686), .C1(new_n676), .C2(new_n681), .ZN(G1330gat));
  OAI211_X1 g486(.A(new_n420), .B(new_n679), .C1(new_n657), .C2(new_n658), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G50gat), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n641), .A2(G50gat), .A3(new_n421), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(KEYINPUT48), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(KEYINPUT105), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n693), .A3(G50gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n691), .B1(new_n698), .B2(new_n699), .ZN(G1331gat));
  AOI21_X1  g499(.A(new_n590), .B1(new_n655), .B2(new_n656), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n663), .A2(new_n613), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(KEYINPUT107), .A3(new_n702), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n643), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n381), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT49), .B(G64gat), .Z(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(G1333gat));
  NAND3_X1  g512(.A1(new_n707), .A2(new_n435), .A3(new_n456), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n705), .A2(new_n628), .A3(new_n706), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G71gat), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n714), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n707), .A2(new_n420), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(G78gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1335gat));
  OAI211_X1 g522(.A(new_n637), .B(new_n702), .C1(new_n657), .C2(new_n658), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(new_n543), .A3(new_n461), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n653), .A2(new_n637), .A3(new_n635), .A4(new_n664), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n614), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n643), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n725), .B1(new_n730), .B2(new_n543), .ZN(G1336gat));
  OAI21_X1  g530(.A(G92gat), .B1(new_n724), .B2(new_n620), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n620), .A2(G92gat), .A3(new_n613), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT52), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n728), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(G1337gat));
  AOI21_X1  g540(.A(G99gat), .B1(new_n729), .B2(new_n456), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n629), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(G99gat), .B2(new_n743), .ZN(G1338gat));
  NOR2_X1   g543(.A1(new_n421), .A2(G106gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G106gat), .B1(new_n724), .B2(new_n421), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT53), .B1(new_n747), .B2(KEYINPUT110), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n748), .B(new_n749), .Z(G1339gat));
  NOR2_X1   g549(.A1(new_n381), .A2(new_n461), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n591), .A2(new_n594), .A3(new_n597), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n599), .A2(KEYINPUT54), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n757));
  AOI21_X1  g556(.A(KEYINPUT97), .B1(new_n595), .B2(new_n598), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n609), .B(new_n597), .C1(new_n591), .C2(new_n594), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n605), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT112), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n763), .A3(new_n605), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n753), .B(new_n756), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n752), .B1(new_n765), .B2(new_n608), .ZN(new_n766));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n760), .B2(new_n605), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n755), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT113), .B(new_n607), .C1(new_n769), .C2(new_n753), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n753), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n766), .A2(new_n663), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n523), .A2(new_n524), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n511), .B1(new_n521), .B2(new_n510), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n530), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n535), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n614), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n635), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n766), .A2(new_n770), .A3(new_n771), .A4(new_n776), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n570), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n637), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n615), .A2(new_n664), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT114), .B1(new_n783), .B2(new_n421), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n785), .B(new_n420), .C1(new_n781), .C2(new_n782), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n456), .B(new_n751), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G113gat), .B1(new_n787), .B2(new_n639), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n751), .ZN(new_n789));
  INV_X1    g588(.A(new_n467), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(G113gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n792), .A3(new_n663), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(G1340gat));
  OAI21_X1  g593(.A(G120gat), .B1(new_n787), .B2(new_n613), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n336), .A3(new_n614), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT115), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n791), .B2(new_n589), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n787), .A2(new_n637), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(G127gat), .ZN(G1342gat));
  NOR4_X1   g600(.A1(new_n789), .A2(G134gat), .A3(new_n790), .A4(new_n570), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT56), .ZN(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n787), .B2(new_n570), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n776), .A2(new_n807), .A3(new_n614), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n535), .A2(new_n775), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n809), .B2(new_n613), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n771), .A2(new_n536), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n607), .B1(new_n769), .B2(new_n753), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n816), .B2(new_n635), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n779), .A2(new_n570), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n812), .A2(new_n814), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n570), .B(new_n819), .C1(new_n820), .C2(new_n811), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n822), .A2(new_n637), .B1(new_n615), .B2(new_n664), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT57), .B1(new_n823), .B2(new_n421), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n783), .A2(new_n825), .A3(new_n420), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n628), .A2(new_n461), .A3(new_n381), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n824), .A2(new_n663), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G141gat), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n628), .A2(new_n421), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT118), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n639), .A2(G141gat), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n783), .A2(new_n751), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n806), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n806), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n824), .A2(new_n536), .A3(new_n826), .A4(new_n827), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(G141gat), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT120), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n839), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n833), .B(KEYINPUT119), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(G141gat), .B2(new_n828), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n841), .B(new_n842), .C1(new_n844), .C2(new_n806), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(G1344gat));
  AND3_X1   g645(.A1(new_n783), .A2(new_n751), .A3(new_n831), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n318), .A3(new_n614), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT121), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n570), .B1(new_n820), .B2(new_n811), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n818), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n818), .B2(new_n852), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n589), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n590), .A2(new_n536), .A3(new_n614), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n825), .B(new_n420), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n783), .A2(new_n420), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n857), .A2(new_n614), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n827), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n850), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT59), .B(new_n318), .C1(new_n863), .C2(new_n614), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n849), .B1(new_n862), .B2(new_n864), .ZN(G1345gat));
  AOI21_X1  g664(.A(G155gat), .B1(new_n847), .B2(new_n589), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n589), .A2(G155gat), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT123), .Z(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n863), .B2(new_n868), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n847), .B2(new_n635), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n863), .A2(G162gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n635), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n643), .B1(new_n781), .B2(new_n782), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n467), .A3(new_n381), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n264), .A3(new_n663), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n784), .A2(new_n786), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n381), .A2(new_n461), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n677), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n536), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(new_n249), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n874), .B2(new_n614), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n614), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT60), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n677), .A2(new_n877), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n784), .B2(new_n786), .ZN(new_n889));
  OAI21_X1  g688(.A(G183gat), .B1(new_n889), .B2(new_n637), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n220), .A3(new_n589), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n886), .A2(KEYINPUT60), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n219), .A3(new_n635), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n635), .B(new_n888), .C1(new_n784), .C2(new_n786), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(G190gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n896), .B2(G190gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT125), .B(new_n895), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1351gat));
  XOR2_X1   g703(.A(KEYINPUT126), .B(G197gat), .Z(new_n905));
  NOR2_X1   g704(.A1(new_n628), .A2(new_n877), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n857), .A2(new_n859), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n639), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n873), .A2(new_n381), .A3(new_n830), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n664), .A2(new_n905), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1352gat));
  AOI21_X1  g711(.A(new_n604), .B1(new_n860), .B2(new_n906), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n604), .A3(new_n614), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT62), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n913), .A2(new_n915), .ZN(G1353gat));
  INV_X1    g715(.A(G211gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n909), .A2(new_n917), .A3(new_n589), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n857), .A2(new_n589), .A3(new_n859), .A4(new_n906), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n909), .B2(new_n635), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n857), .A2(new_n924), .A3(new_n859), .A4(new_n906), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n205), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n570), .B1(new_n907), .B2(KEYINPUT127), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1355gat));
endmodule


