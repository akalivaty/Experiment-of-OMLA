//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n193), .A2(new_n206), .A3(new_n209), .A4(new_n197), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G134), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(new_n214), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n218), .B2(G134), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n215), .A3(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n215), .A2(G137), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n224), .A2(new_n226), .B1(new_n227), .B2(KEYINPUT11), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n222), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n223), .B1(new_n222), .B2(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT12), .B1(new_n213), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n229), .B2(new_n230), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT12), .B1(new_n211), .B2(new_n212), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n220), .B1(new_n219), .B2(new_n214), .ZN(new_n236));
  AOI211_X1 g050(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n218), .C2(G134), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n226), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n227), .A2(KEYINPUT11), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n222), .A2(new_n223), .A3(new_n228), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT68), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n232), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n234), .A2(new_n244), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT0), .A4(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n190), .A2(new_n192), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G128), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n257), .A3(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n210), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n193), .A2(new_n197), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT10), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n263));
  NAND2_X1  g077(.A1(new_n212), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n248), .A2(KEYINPUT83), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n234), .A2(new_n244), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n247), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT81), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n268), .A2(new_n269), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT83), .B1(new_n248), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(new_n267), .A3(new_n269), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n187), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  INV_X1    g102(.A(new_n279), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n266), .B2(new_n270), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n277), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n247), .B(new_n276), .C1(new_n266), .C2(new_n270), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT84), .B(G469), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n292), .B1(new_n276), .B2(new_n282), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n288), .A3(new_n285), .A4(new_n295), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G221), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n285), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(KEYINPUT86), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n280), .A2(new_n281), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n276), .B1(new_n308), .B2(new_n289), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n277), .B(new_n246), .C1(new_n280), .C2(new_n281), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n285), .B(new_n295), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT85), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n286), .B1(new_n312), .B2(new_n298), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n313), .B2(new_n304), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G210), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G119), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT67), .B1(new_n322), .B2(G116), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n320), .A3(G119), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n327));
  INV_X1    g141(.A(G113), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n321), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT2), .B(G113), .Z(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n260), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n326), .A2(new_n332), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n326), .A2(new_n332), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n258), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n251), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n255), .A2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n261), .B2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n274), .A2(G224), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n339), .A2(KEYINPUT87), .A3(new_n341), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n334), .B(new_n340), .C1(new_n337), .C2(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT6), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT87), .B1(new_n339), .B2(new_n341), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT88), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n349), .A2(KEYINPUT6), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(new_n348), .ZN(new_n356));
  AOI211_X1 g170(.A(new_n343), .B(new_n347), .C1(new_n352), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(KEYINPUT7), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n345), .B(new_n358), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n340), .B(KEYINPUT8), .ZN(new_n360));
  INV_X1    g174(.A(new_n334), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n260), .B1(new_n331), .B2(new_n333), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n363), .A3(new_n349), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n285), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n319), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n352), .A2(new_n356), .ZN(new_n367));
  INV_X1    g181(.A(new_n343), .ZN(new_n368));
  INV_X1    g182(.A(new_n347), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n365), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n318), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n317), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G475), .ZN(new_n374));
  XNOR2_X1  g188(.A(G125), .B(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n191), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(KEYINPUT79), .Z(new_n377));
  INV_X1    g191(.A(G125), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n378), .A2(KEYINPUT77), .A3(G140), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G146), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n274), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n188), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n384), .A2(new_n274), .A3(G143), .A4(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  OR3_X1    g203(.A1(new_n388), .A2(KEYINPUT89), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n388), .B2(KEYINPUT89), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G125), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT78), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n378), .A2(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n395), .A3(new_n380), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n378), .A2(KEYINPUT77), .A3(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n400), .B2(KEYINPUT16), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT16), .ZN(new_n402));
  AOI211_X1 g216(.A(KEYINPUT78), .B(new_n402), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  OAI21_X1  g217(.A(G146), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n396), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n381), .B2(new_n402), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT78), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n191), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n388), .A2(KEYINPUT17), .A3(G131), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n388), .A2(G131), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n386), .A2(new_n223), .A3(new_n387), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n404), .A2(new_n409), .A3(new_n410), .A4(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n199), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n393), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n393), .B2(new_n415), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n374), .B1(new_n421), .B2(new_n285), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n191), .B1(new_n406), .B2(new_n408), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n375), .A2(KEYINPUT19), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n400), .B2(KEYINPUT19), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G146), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT91), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n425), .A2(G146), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n404), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n411), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT90), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n411), .A2(new_n433), .A3(new_n413), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n417), .B1(new_n436), .B2(new_n393), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n419), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT20), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n439), .C1(new_n437), .C2(new_n419), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n422), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G952), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  INV_X1    g260(.A(G234), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(new_n384), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G898), .Z(new_n449));
  OAI211_X1 g263(.A(G902), .B(G953), .C1(new_n447), .C2(new_n384), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT92), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n320), .A2(G122), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n455), .B2(KEYINPUT14), .ZN(new_n458));
  OR3_X1    g272(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT14), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(new_n456), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G107), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n202), .A3(new_n455), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT93), .ZN(new_n463));
  XNOR2_X1  g277(.A(G128), .B(G143), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n215), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n454), .A2(new_n466), .A3(new_n202), .A4(new_n455), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n461), .A2(new_n463), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT13), .B1(new_n196), .B2(G143), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n215), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n464), .ZN(new_n471));
  INV_X1    g285(.A(new_n462), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n202), .B1(new_n454), .B2(new_n455), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n303), .A2(G217), .A3(new_n274), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n285), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n486), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(new_n285), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n444), .A2(new_n451), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n373), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT96), .B1(new_n315), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G217), .B1(new_n447), .B2(G902), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT74), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n322), .A2(G128), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT23), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT75), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n322), .A2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT76), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT76), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n502), .A2(new_n322), .A3(G128), .ZN(new_n510));
  OAI21_X1  g324(.A(G110), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT24), .B(G110), .Z(new_n512));
  XNOR2_X1  g326(.A(G119), .B(G128), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n401), .A2(new_n403), .A3(G146), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n511), .B(new_n514), .C1(new_n515), .C2(new_n423), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n509), .A2(G110), .A3(new_n510), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n512), .A2(new_n513), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n404), .B(new_n377), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n301), .A2(new_n447), .A3(G953), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  AND3_X1   g336(.A1(new_n516), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n516), .B2(new_n519), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT25), .B1(new_n525), .B2(new_n285), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(new_n519), .ZN(new_n527));
  INV_X1    g341(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n519), .A3(new_n522), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n498), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT80), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n285), .A3(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n531), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n498), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n498), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n525), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n326), .B(new_n332), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n256), .B1(new_n229), .B2(new_n230), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT66), .ZN(new_n547));
  XNOR2_X1  g361(.A(G134), .B(G137), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n223), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n218), .A2(G134), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT66), .B(G131), .C1(new_n227), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n261), .A2(new_n243), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n234), .A2(new_n256), .A3(new_n244), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n261), .A2(new_n243), .A3(new_n552), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n544), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n556), .A2(new_n560), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n384), .A2(new_n274), .A3(G210), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT27), .Z(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT69), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n557), .A2(new_n561), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n557), .A2(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n255), .B1(new_n242), .B2(new_n243), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n555), .B1(new_n571), .B2(new_n558), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n544), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n569), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n566), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n557), .A2(new_n561), .B1(new_n554), .B2(new_n544), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n579), .B(new_n567), .C1(new_n580), .C2(new_n578), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT70), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT70), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n576), .A4(new_n568), .ZN(new_n587));
  INV_X1    g401(.A(new_n569), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n545), .B1(new_n557), .B2(new_n553), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT28), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n569), .A2(KEYINPUT71), .A3(new_n578), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n566), .A2(new_n582), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n285), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n584), .A2(new_n587), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT72), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n601), .A3(G472), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n567), .B(new_n569), .C1(new_n570), .C2(new_n573), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT31), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n562), .A2(KEYINPUT31), .A3(new_n567), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n579), .B1(new_n580), .B2(new_n578), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n566), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(G472), .A2(G902), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(KEYINPUT32), .A3(new_n612), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT32), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n606), .A2(new_n607), .B1(new_n566), .B2(new_n609), .ZN(new_n616));
  INV_X1    g430(.A(new_n612), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n619), .B2(KEYINPUT73), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n543), .B1(new_n603), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n315), .A2(KEYINPUT96), .A3(new_n494), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n496), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NOR3_X1   g438(.A1(new_n357), .A2(new_n365), .A3(new_n319), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n318), .B1(new_n370), .B2(new_n371), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n316), .B(new_n451), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n480), .B(KEYINPUT33), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n482), .A2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(G478), .B1(new_n480), .B2(new_n285), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n421), .A2(new_n285), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G475), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n432), .A2(new_n434), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n428), .A2(new_n404), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n639), .B2(KEYINPUT91), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n640), .A2(new_n430), .B1(new_n383), .B2(new_n392), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n418), .B1(new_n641), .B2(new_n417), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n442), .B1(new_n642), .B2(new_n439), .ZN(new_n643));
  INV_X1    g457(.A(new_n443), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n627), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n616), .B2(G902), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n616), .B2(new_n617), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n543), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n315), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n642), .A2(new_n654), .A3(new_n442), .A4(new_n439), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n443), .A2(KEYINPUT98), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n441), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n656), .A3(new_n441), .A4(KEYINPUT99), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n637), .A2(new_n490), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n627), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n315), .A2(new_n665), .A3(new_n650), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n539), .B1(new_n538), .B2(new_n498), .ZN(new_n670));
  INV_X1    g484(.A(new_n498), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT80), .B(new_n671), .C1(new_n537), .C2(new_n531), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n527), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n541), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n669), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n534), .A2(new_n669), .A3(new_n540), .A4(new_n676), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n677), .A2(new_n679), .A3(new_n649), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n496), .A2(new_n622), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NAND2_X1  g497(.A1(new_n366), .A2(new_n372), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n316), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n677), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(G472), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n568), .A2(new_n576), .A3(new_n582), .A4(new_n581), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n596), .B1(new_n688), .B2(KEYINPUT70), .ZN(new_n689));
  AOI211_X1 g503(.A(KEYINPUT72), .B(new_n687), .C1(new_n689), .C2(new_n587), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n601), .B1(new_n598), .B2(G472), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n620), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n448), .B(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(G900), .B2(new_n450), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT102), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n664), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n686), .A2(new_n692), .A3(new_n315), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n695), .B(KEYINPUT39), .Z(new_n699));
  AND2_X1   g513(.A1(new_n315), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n588), .A2(new_n589), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n604), .B1(new_n703), .B2(new_n567), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n285), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n620), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n684), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n534), .A2(new_n540), .A3(new_n676), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n444), .A2(new_n491), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n316), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n708), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n700), .A2(new_n701), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n702), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  INV_X1    g532(.A(new_n695), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n635), .A2(new_n645), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n686), .A2(new_n692), .A3(new_n315), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT104), .B(G146), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G48));
  NAND2_X1  g538(.A1(new_n312), .A2(new_n298), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n293), .A2(new_n187), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n305), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n543), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n692), .A2(new_n647), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n692), .A2(new_n731), .A3(new_n647), .A4(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT106), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n733), .B(new_n735), .ZN(G15));
  NAND3_X1  g550(.A1(new_n692), .A2(new_n665), .A3(new_n728), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  NAND2_X1  g552(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n492), .A3(new_n678), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n685), .A2(new_n727), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n692), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n373), .A2(new_n713), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n725), .A2(new_n305), .A3(new_n451), .A4(new_n726), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n567), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n608), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n612), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n648), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n673), .A2(KEYINPUT108), .A3(new_n542), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n543), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n746), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NOR2_X1   g574(.A1(new_n753), .A2(new_n712), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n721), .A3(new_n741), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  AOI21_X1  g577(.A(new_n246), .B1(new_n280), .B2(new_n281), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT109), .B1(new_n764), .B2(new_n276), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n271), .A2(new_n766), .A3(new_n277), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n767), .A3(new_n283), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n285), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(G469), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n304), .B1(new_n725), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n366), .A2(new_n316), .A3(new_n372), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n721), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n619), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n690), .B2(new_n691), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n776), .A3(new_n758), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n773), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(KEYINPUT42), .A3(new_n720), .ZN(new_n779));
  AOI22_X1  g593(.A1(KEYINPUT42), .A2(new_n777), .B1(new_n621), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  INV_X1    g595(.A(new_n778), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n696), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT110), .B1(new_n664), .B2(new_n695), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n621), .A2(new_n782), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n187), .B1(new_n284), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n788), .B2(new_n768), .ZN(new_n790));
  NAND2_X1  g604(.A1(G469), .A2(G902), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n725), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n305), .B(new_n699), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n796), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n802), .B2(new_n794), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n305), .A4(new_n699), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n635), .A2(new_n444), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT43), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n649), .A3(new_n711), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n811), .A2(new_n812), .A3(new_n772), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  INV_X1    g629(.A(new_n543), .ZN(new_n816));
  OR4_X1    g630(.A1(new_n692), .A2(new_n816), .A3(new_n720), .A4(new_n772), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n803), .B2(new_n304), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT47), .B(new_n305), .C1(new_n797), .C2(new_n798), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(new_n394), .ZN(G42));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n730), .A2(new_n732), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n742), .A2(new_n737), .A3(new_n759), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n742), .A2(new_n737), .A3(new_n759), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n733), .A2(new_n827), .A3(KEYINPUT113), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n777), .A2(KEYINPUT42), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n621), .A2(new_n779), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n786), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n627), .B2(new_n646), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n645), .A2(new_n491), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n373), .A2(new_n451), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n635), .A2(new_n645), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n373), .A3(KEYINPUT114), .A4(new_n451), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n839), .A2(new_n315), .A3(new_n650), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n315), .A2(KEYINPUT96), .A3(new_n494), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n495), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n842), .B2(new_n621), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n677), .A2(new_n679), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n490), .A2(new_n422), .A3(new_n695), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n366), .A2(new_n845), .A3(new_n372), .A4(new_n316), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n659), .B2(new_n660), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n692), .A2(new_n315), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n846), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n661), .A2(new_n851), .A3(new_n739), .A4(new_n678), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .A3(new_n692), .A4(new_n315), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n850), .A2(new_n853), .B1(new_n761), .B2(new_n774), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n832), .A2(new_n843), .A3(new_n854), .A4(new_n681), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT116), .B1(new_n829), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n733), .A2(new_n827), .A3(KEYINPUT113), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT113), .B1(new_n733), .B2(new_n827), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n853), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n774), .A2(new_n761), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n780), .A3(new_n786), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n840), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n623), .A2(new_n681), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n744), .A2(new_n711), .A3(new_n695), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n707), .A3(new_n771), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n697), .A2(new_n722), .A3(new_n762), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(KEYINPUT117), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n856), .A2(new_n867), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n856), .A2(new_n867), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n881), .B(KEYINPUT54), .C1(new_n882), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n884), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n824), .A2(new_n825), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n865), .A2(new_n883), .A3(KEYINPUT53), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(KEYINPUT54), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n693), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n808), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n727), .A2(new_n772), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n893), .A2(new_n761), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n543), .A2(new_n448), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n708), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(new_n645), .A3(new_n635), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n725), .A2(new_n726), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n819), .B(new_n820), .C1(new_n305), .C2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n754), .A3(new_n758), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n772), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n895), .B(new_n898), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n316), .B1(KEYINPUT118), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n710), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n901), .A2(new_n727), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n903), .A2(KEYINPUT51), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n893), .A2(new_n758), .A3(new_n776), .A4(new_n894), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT48), .Z(new_n912));
  INV_X1    g726(.A(new_n741), .ZN(new_n913));
  OAI221_X1 g727(.A(new_n446), .B1(new_n646), .B2(new_n897), .C1(new_n901), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n909), .B(KEYINPUT119), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n903), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n910), .B(new_n915), .C1(new_n917), .C2(KEYINPUT51), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n891), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n807), .A2(new_n304), .A3(new_n317), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n710), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n899), .A2(KEYINPUT49), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n755), .A2(new_n757), .B1(KEYINPUT49), .B2(new_n899), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n921), .A2(new_n708), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G75));
  NAND2_X1  g739(.A1(new_n445), .A2(G953), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT121), .Z(new_n927));
  AOI21_X1  g741(.A(new_n285), .B1(new_n887), .B2(new_n889), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n343), .B1(new_n352), .B2(new_n356), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n369), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n357), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n927), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n928), .A2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n929), .A2(KEYINPUT120), .A3(new_n933), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G51));
  INV_X1    g755(.A(new_n927), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n791), .B(KEYINPUT57), .Z(new_n943));
  NOR2_X1   g757(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n944));
  INV_X1    g758(.A(new_n889), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n880), .B2(new_n884), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n297), .ZN(new_n950));
  INV_X1    g764(.A(new_n928), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(new_n790), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n942), .B1(new_n950), .B2(new_n952), .ZN(G54));
  NAND2_X1  g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n642), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .A4(new_n438), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n942), .B1(new_n955), .B2(new_n956), .ZN(G60));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n628), .B(new_n960), .C1(new_n944), .C2(new_n948), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n927), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n628), .B1(new_n891), .B2(new_n960), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n946), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(new_n525), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n942), .B1(new_n967), .B2(new_n675), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT122), .B1(new_n967), .B2(new_n675), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(KEYINPUT61), .ZN(new_n971));
  INV_X1    g785(.A(new_n966), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n890), .A2(new_n675), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n973), .B(new_n927), .C1(new_n525), .C2(new_n967), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT61), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n977), .ZN(G66));
  AOI21_X1  g792(.A(new_n274), .B1(new_n449), .B2(G224), .ZN(new_n979));
  INV_X1    g793(.A(new_n864), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n859), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(new_n274), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n930), .B1(new_n983), .B2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n560), .A2(new_n572), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n425), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n821), .B1(new_n806), .B2(new_n813), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n697), .A2(new_n762), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n722), .ZN(new_n991));
  AND4_X1   g805(.A1(new_n373), .A2(new_n776), .A3(new_n713), .A4(new_n758), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n806), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n832), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n989), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n987), .B(new_n988), .C1(new_n997), .C2(G953), .ZN(new_n998));
  INV_X1    g812(.A(new_n835), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n772), .B1(new_n999), .B2(new_n646), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n700), .A2(new_n621), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n991), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n717), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n989), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(G953), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n998), .B1(new_n1010), .B2(new_n987), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1012), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1014), .B(new_n998), .C1(new_n1010), .C2(new_n987), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G72));
  XNOR2_X1  g830(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n687), .A2(new_n285), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1017), .B(new_n1018), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n997), .B2(new_n981), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n562), .B(KEYINPUT126), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n566), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1019), .ZN(new_n1024));
  INV_X1    g838(.A(new_n981), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1009), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1021), .A2(new_n567), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n927), .B(new_n1023), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n882), .A2(new_n885), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(KEYINPUT53), .B2(new_n880), .ZN(new_n1030));
  INV_X1    g844(.A(new_n577), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1024), .B1(new_n1031), .B2(new_n604), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(G57));
endmodule


