//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n192), .A2(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(G143), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n197), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n196), .A2(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n204), .A3(G128), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n189), .A2(new_n191), .B1(new_n188), .B2(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n212));
  INV_X1    g026(.A(G224), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G953), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT85), .A3(G224), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n211), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G104), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(G107), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(G104), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n219), .A2(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT2), .B(G113), .Z(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT5), .ZN(new_n238));
  OR3_X1    g052(.A1(new_n235), .A2(KEYINPUT5), .A3(G119), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g056(.A(G110), .B(G122), .Z(new_n243));
  XOR2_X1   g057(.A(new_n243), .B(KEYINPUT8), .Z(new_n244));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT82), .A4(G113), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n237), .A3(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n242), .B(new_n244), .C1(new_n248), .C2(new_n231), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n220), .A2(new_n223), .A3(new_n225), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n220), .A2(new_n223), .A3(KEYINPUT78), .A4(new_n225), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(G101), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n252), .A2(KEYINPUT4), .A3(G101), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n234), .A2(new_n236), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT2), .B(G113), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n237), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n237), .A2(KEYINPUT68), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n248), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n226), .A2(new_n229), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n226), .B2(new_n229), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n258), .A2(new_n266), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n243), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT83), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n256), .A2(new_n257), .B1(new_n264), .B2(new_n265), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n269), .A2(new_n270), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n248), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  NOR4_X1   g092(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n243), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n218), .B(new_n249), .C1(new_n274), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n258), .A2(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n267), .A2(new_n271), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(new_n243), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n274), .B2(new_n279), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n283), .A3(new_n243), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n214), .A2(new_n216), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n290), .B(KEYINPUT84), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n211), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT86), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(new_n296), .A3(new_n289), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n282), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT88), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n282), .ZN(new_n301));
  INV_X1    g115(.A(new_n289), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n284), .A2(new_n273), .A3(new_n285), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n278), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n272), .A2(KEYINPUT83), .A3(new_n273), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n306), .B2(new_n287), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n307), .B2(new_n293), .ZN(new_n308));
  INV_X1    g122(.A(new_n297), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n301), .B(new_n299), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n299), .B(KEYINPUT87), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n298), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n300), .B1(new_n312), .B2(KEYINPUT88), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT96), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(G953), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n188), .A2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n195), .A2(G143), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G134), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n320), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n324), .A2(KEYINPUT93), .A3(G134), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT13), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n320), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n319), .A2(new_n327), .ZN(new_n330));
  OAI21_X1  g144(.A(G134), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n332));
  INV_X1    g146(.A(G122), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(G116), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n235), .A2(KEYINPUT92), .A3(G122), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n334), .A2(new_n335), .B1(G116), .B2(new_n333), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(G107), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(G107), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n326), .B(new_n331), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT14), .B1(new_n334), .B2(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n340), .A3(G107), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n324), .B(G134), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n222), .A2(KEYINPUT14), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n341), .B(new_n342), .C1(new_n336), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n317), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n339), .A2(new_n344), .A3(new_n317), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AND4_X1   g163(.A1(KEYINPUT94), .A2(new_n339), .A3(new_n344), .A4(new_n317), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n351), .A3(new_n281), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT95), .A4(new_n281), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G478), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT15), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n352), .A2(new_n358), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n215), .A3(G214), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n188), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n369), .B2(KEYINPUT16), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT16), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(new_n368), .A3(KEYINPUT75), .A4(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n209), .A2(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n370), .B(new_n372), .C1(new_n374), .C2(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n190), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n369), .A2(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(G146), .A3(new_n370), .A4(new_n372), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n366), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n366), .A2(new_n376), .A3(new_n379), .A4(KEYINPUT91), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n365), .A2(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n364), .B(G143), .ZN(new_n385));
  INV_X1    g199(.A(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n382), .B(new_n383), .C1(KEYINPUT17), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n219), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n385), .B1(new_n392), .B2(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n377), .A2(new_n190), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n374), .A2(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n393), .B(new_n396), .C1(new_n392), .C2(new_n384), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n391), .B1(new_n389), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n281), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G475), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT21), .B(G898), .Z(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G234), .A2(G237), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(G902), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n215), .A2(G952), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n404), .A2(new_n407), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n377), .A2(KEYINPUT90), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT19), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n388), .A2(new_n379), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n397), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n391), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G475), .B1(new_n398), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(new_n281), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n418), .B2(new_n281), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n402), .B(new_n410), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n314), .B1(new_n362), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n281), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n419), .A3(new_n281), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n427), .A2(new_n428), .B1(G475), .B2(new_n401), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n360), .B1(new_n356), .B2(new_n358), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT96), .A4(new_n410), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n313), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT24), .B(G110), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G119), .B(G128), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n376), .A2(new_n379), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n233), .A2(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT23), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT74), .B1(new_n195), .B2(G119), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G110), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n438), .A2(new_n439), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n444), .A2(G110), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n379), .B(new_n394), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT22), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(G137), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n449), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n281), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT25), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n316), .B1(G234), .B2(new_n281), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT25), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n455), .A2(new_n456), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n462), .A2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT77), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT11), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n322), .B2(G137), .ZN(new_n473));
  INV_X1    g287(.A(G137), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT11), .A3(G134), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n322), .A2(G137), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n386), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n474), .A2(G134), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n322), .A2(G137), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n477), .B2(new_n480), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n476), .A3(new_n475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G131), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n477), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n484), .A2(new_n208), .B1(new_n202), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n471), .B1(new_n488), .B2(KEYINPUT30), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n196), .A2(new_n198), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n200), .A2(new_n201), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n202), .A2(KEYINPUT69), .A3(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n208), .A2(new_n477), .A3(new_n480), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT30), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n477), .A2(new_n480), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT66), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n208), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n492), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(KEYINPUT67), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n489), .A2(new_n266), .A3(new_n497), .A4(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n266), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n494), .A3(new_n496), .A4(new_n495), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n363), .A2(new_n215), .A3(G210), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT27), .Z(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT26), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n224), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n508), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(KEYINPUT70), .A3(new_n507), .A4(new_n512), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n502), .A2(new_n266), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT28), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n496), .A2(new_n492), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT28), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n512), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n513), .A2(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G472), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n281), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n470), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n514), .A2(new_n515), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n514), .A2(new_n515), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(KEYINPUT32), .A3(new_n526), .A4(new_n281), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n508), .A2(new_n512), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n523), .A2(new_n524), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT29), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n266), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n507), .ZN(new_n540));
  OR3_X1    g354(.A1(new_n537), .A2(new_n539), .A3(new_n266), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n522), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n512), .A2(KEYINPUT29), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n281), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G472), .B1(new_n536), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n528), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT72), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n528), .A2(new_n533), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n469), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT79), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n195), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n555), .B2(new_n554), .ZN(new_n557));
  INV_X1    g371(.A(new_n200), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n230), .B1(new_n559), .B2(new_n205), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT10), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n258), .A2(new_n202), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n208), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n487), .B(KEYINPUT81), .Z(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n487), .B1(new_n567), .B2(new_n561), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  INV_X1    g383(.A(G227), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n569), .B(new_n571), .Z(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n567), .A2(new_n561), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n208), .A2(new_n231), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n487), .B1(new_n560), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT12), .B(new_n487), .C1(new_n560), .C2(new_n575), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n574), .A2(new_n565), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n573), .B(G469), .C1(new_n580), .C2(new_n572), .ZN(new_n581));
  NAND2_X1  g395(.A1(G469), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G469), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n566), .A3(new_n572), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n572), .B1(new_n566), .B2(new_n568), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n585), .B(new_n281), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n553), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n435), .A2(new_n551), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NAND2_X1  g407(.A1(new_n356), .A2(new_n357), .ZN(new_n594));
  INV_X1    g408(.A(new_n348), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n346), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n348), .A2(KEYINPUT98), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT33), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT33), .B1(new_n349), .B2(new_n351), .ZN(new_n601));
  OAI211_X1 g415(.A(G478), .B(new_n281), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n402), .B1(new_n420), .B2(new_n423), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n603), .A2(KEYINPUT99), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT99), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT97), .B1(new_n298), .B2(new_n299), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n610));
  INV_X1    g424(.A(new_n299), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n310), .ZN(new_n613));
  AND4_X1   g427(.A1(new_n433), .A2(new_n607), .A3(new_n613), .A4(new_n410), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n525), .B2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n532), .A2(new_n526), .A3(new_n281), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n469), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n617), .A2(new_n618), .A3(new_n591), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  XNOR2_X1  g436(.A(new_n426), .B(new_n421), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n402), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n430), .ZN(new_n625));
  AND4_X1   g439(.A1(new_n433), .A2(new_n613), .A3(new_n410), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n619), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n454), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n450), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n467), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n464), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(KEYINPUT100), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(KEYINPUT100), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n435), .A2(new_n591), .A3(new_n617), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT37), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(G110), .Z(G12));
  AOI21_X1  g454(.A(new_n636), .B1(new_n548), .B2(new_n550), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n613), .A2(new_n433), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n408), .A2(new_n405), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT101), .Z(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n407), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n624), .A2(new_n430), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(new_n591), .A3(new_n642), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XNOR2_X1  g463(.A(new_n313), .B(KEYINPUT38), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(G902), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n505), .A2(new_n507), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n512), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n528), .A2(new_n533), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n650), .A2(new_n633), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n646), .B(KEYINPUT39), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n591), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n429), .A2(new_n430), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n434), .B1(new_n662), .B2(KEYINPUT40), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n659), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  INV_X1    g482(.A(new_n646), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n603), .A2(new_n604), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n642), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n613), .A2(new_n433), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT102), .B1(new_n673), .B2(new_n670), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n591), .A3(new_n674), .A4(new_n641), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  NOR2_X1   g490(.A1(new_n588), .A2(new_n589), .ZN(new_n677));
  OAI21_X1  g491(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n552), .A3(new_n590), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n614), .A2(new_n551), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NAND3_X1  g496(.A1(new_n626), .A2(new_n551), .A3(new_n679), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT103), .B(G116), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G18));
  INV_X1    g499(.A(new_n432), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n613), .A2(new_n433), .A3(new_n679), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n641), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  AND3_X1   g503(.A1(new_n613), .A2(new_n433), .A3(new_n664), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n513), .A2(new_n516), .B1(new_n543), .B2(new_n524), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(new_n527), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n615), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n618), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n690), .A2(new_n694), .A3(new_n410), .A4(new_n679), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  AND3_X1   g510(.A1(new_n693), .A2(new_n633), .A3(new_n671), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n687), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  NAND2_X1  g513(.A1(new_n295), .A2(new_n297), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n311), .B1(new_n700), .B2(new_n301), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n611), .B(new_n282), .C1(new_n295), .C2(new_n297), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT88), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n300), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n584), .A2(KEYINPUT104), .A3(new_n590), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n566), .A2(new_n568), .ZN(new_n707));
  INV_X1    g521(.A(new_n572), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(G469), .B(G902), .C1(new_n709), .C2(new_n587), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n706), .B1(new_n710), .B2(new_n583), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n553), .A2(new_n434), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n703), .A2(new_n704), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n313), .A2(KEYINPUT105), .A3(new_n712), .A4(new_n713), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n551), .A3(new_n671), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n547), .A2(new_n618), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n670), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n722), .A2(new_n718), .A3(KEYINPUT42), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n720), .B1(new_n716), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n721), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NAND3_X1  g543(.A1(new_n718), .A2(new_n551), .A3(new_n647), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  INV_X1    g545(.A(KEYINPUT33), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n595), .A2(new_n345), .A3(KEYINPUT94), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n350), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n357), .B(G902), .C1(new_n734), .C2(new_n599), .ZN(new_n735));
  AOI21_X1  g549(.A(G478), .B1(new_n354), .B2(new_n355), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n604), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n615), .A2(new_n616), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n633), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT108), .Z(new_n744));
  OAI21_X1  g558(.A(new_n573), .B1(new_n580), .B2(new_n572), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n747), .B2(new_n582), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n710), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n582), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n552), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n660), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n313), .A2(new_n433), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n741), .B2(new_n742), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n744), .A2(new_n753), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND3_X1  g574(.A1(new_n548), .A2(new_n550), .A3(new_n671), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n618), .A3(new_n754), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT110), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  AND4_X1   g582(.A1(new_n618), .A2(new_n658), .A3(new_n713), .A4(new_n738), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n678), .A2(new_n590), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT49), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n650), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n718), .A2(new_n697), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n591), .A2(new_n402), .A3(new_n623), .A4(new_n669), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n641), .A2(new_n755), .A3(new_n430), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n680), .A2(new_n683), .A3(new_n688), .A4(new_n695), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n604), .A2(new_n430), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT111), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n429), .B2(new_n737), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n313), .A2(new_n434), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n619), .A3(new_n782), .A4(new_n410), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n638), .A2(new_n592), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n728), .A2(new_n730), .A3(new_n777), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n658), .A2(new_n633), .A3(new_n646), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n690), .A3(new_n552), .A4(new_n712), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n675), .A2(new_n648), .A3(new_n698), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n778), .A2(new_n776), .A3(new_n784), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n795), .A3(new_n728), .A4(new_n730), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n791), .B2(new_n792), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(KEYINPUT113), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n787), .A4(new_n796), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n797), .A2(new_n805), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n728), .A2(new_n730), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n810), .A4(new_n794), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n694), .A2(new_n644), .A3(new_n739), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n650), .A3(new_n434), .A4(new_n679), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT50), .Z(new_n816));
  AND4_X1   g630(.A1(new_n644), .A2(new_n755), .A3(new_n679), .A4(new_n739), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n633), .A3(new_n693), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n755), .A2(new_n618), .A3(new_n679), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n643), .A3(new_n657), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n429), .A3(new_n737), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n770), .A2(new_n553), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n764), .B2(new_n765), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n755), .A3(new_n814), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(KEYINPUT51), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT117), .ZN(new_n829));
  INV_X1    g643(.A(new_n723), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n817), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT48), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n820), .A2(new_n607), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n817), .A2(new_n830), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n833), .A2(new_n408), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n822), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n814), .A2(new_n687), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n828), .A2(KEYINPUT117), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n813), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(G952), .A2(G953), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n772), .B1(new_n847), .B2(new_n848), .ZN(G75));
  AOI21_X1  g663(.A(new_n281), .B1(new_n808), .B2(new_n811), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n850), .B2(G210), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n307), .B(new_n293), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT55), .Z(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n215), .A2(G952), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT119), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n311), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n854), .A2(new_n856), .A3(new_n860), .ZN(G51));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n582), .B(KEYINPUT57), .Z(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n808), .A2(new_n811), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(new_n812), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n867), .B2(new_n677), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n850), .A2(G469), .A3(new_n746), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n677), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n855), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(G54));
  NAND3_X1  g691(.A1(new_n850), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n398), .A2(new_n417), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n878), .A2(new_n880), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n855), .ZN(G60));
  NAND2_X1  g698(.A1(G478), .A2(G902), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT59), .Z(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n600), .A2(new_n601), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n866), .B2(new_n812), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n807), .B2(new_n812), .ZN(new_n890));
  INV_X1    g704(.A(new_n888), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n890), .A2(KEYINPUT122), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT122), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  AOI221_X4 g707(.A(new_n856), .B1(new_n887), .B2(new_n889), .C1(new_n892), .C2(new_n893), .ZN(G63));
  INV_X1    g708(.A(new_n856), .ZN(new_n895));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT60), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n808), .B2(new_n811), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n465), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n631), .B2(new_n898), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g715(.A(G953), .B1(new_n404), .B2(new_n213), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n785), .B2(G953), .ZN(new_n903));
  INV_X1    g717(.A(new_n307), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(G898), .B2(new_n215), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(G69));
  XNOR2_X1  g720(.A(new_n810), .B(KEYINPUT123), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n675), .A2(new_n648), .A3(new_n698), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n766), .A2(new_n759), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n753), .A2(new_n690), .A3(new_n830), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n489), .A2(new_n497), .A3(new_n504), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n412), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n215), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n666), .A2(new_n908), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT62), .Z(new_n916));
  INV_X1    g730(.A(new_n662), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n551), .A2(new_n755), .A3(new_n781), .A4(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n918), .A3(new_n909), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n215), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n913), .B1(G900), .B2(new_n215), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n570), .B2(new_n645), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n914), .A2(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n923), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT125), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G72));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  INV_X1    g744(.A(new_n785), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n911), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n653), .A2(new_n512), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n855), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n930), .B1(new_n919), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n655), .ZN(new_n936));
  INV_X1    g750(.A(new_n930), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n655), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT126), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n798), .A2(new_n806), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G57));
endmodule


