//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OR3_X1    g038(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT68), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n472), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n472), .A2(G138), .ZN(new_n485));
  XOR2_X1   g060(.A(KEYINPUT69), .B(KEYINPUT4), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n472), .B(G138), .C1(KEYINPUT69), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n479), .B2(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT70), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT70), .A2(G543), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n501), .B(KEYINPUT5), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n497), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n500), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT72), .Z(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AND3_X1   g098(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n524));
  AOI211_X1 g099(.A(new_n523), .B(new_n524), .C1(G51), .C2(new_n499), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n512), .A2(new_n497), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n516), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n526), .A2(G90), .B1(G52), .B2(new_n499), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AND2_X1   g108(.A1(new_n512), .A2(G56), .ZN(new_n534));
  AND2_X1   g109(.A1(G68), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n512), .A2(G81), .A3(new_n497), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT73), .B(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n499), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n537), .A2(KEYINPUT74), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT74), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n512), .A2(G91), .A3(new_n497), .ZN(new_n550));
  AND2_X1   g125(.A1(G78), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n512), .B2(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n552), .B2(new_n516), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT75), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n558), .A2(new_n497), .A3(G53), .A4(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT6), .A2(G651), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n555), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n559), .A2(new_n563), .A3(KEYINPUT76), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT76), .B1(new_n559), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n549), .B1(new_n553), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n559), .A2(new_n563), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n559), .A2(new_n563), .A3(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT5), .B1(new_n502), .B2(new_n503), .ZN(new_n574));
  INV_X1    g149(.A(new_n511), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(new_n504), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n577), .B2(new_n551), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n572), .A2(KEYINPUT77), .A3(new_n578), .A4(new_n550), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n567), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n525), .A2(new_n527), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  AND3_X1   g158(.A1(new_n526), .A2(KEYINPUT78), .A3(G87), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n526), .B2(G87), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n512), .A2(G74), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G49), .B2(new_n499), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n526), .A2(G86), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n499), .A2(G48), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n516), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n516), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n526), .A2(G85), .B1(G47), .B2(new_n499), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G301), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n512), .A2(G66), .ZN(new_n603));
  INV_X1    g178(.A(G79), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n507), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n499), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n512), .A2(G92), .A3(new_n497), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT80), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n602), .B1(new_n611), .B2(new_n601), .ZN(G284));
  AOI21_X1  g187(.A(new_n602), .B1(new_n611), .B2(new_n601), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n580), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n580), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n611), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  INV_X1    g198(.A(new_n469), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n473), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n472), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n479), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n478), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT86), .Z(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2451), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n647), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(G14), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n629), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n637), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n674), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n674), .A2(new_n682), .ZN(new_n684));
  NOR4_X1   g259(.A1(new_n680), .A2(new_n681), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1981), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G34), .ZN(new_n692));
  AOI21_X1  g267(.A(G29), .B1(new_n692), .B2(KEYINPUT24), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(KEYINPUT24), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n475), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G11), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT102), .B(G28), .Z(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n701), .B2(KEYINPUT30), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(KEYINPUT30), .B2(new_n701), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n703), .C1(new_n636), .C2(new_n695), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(G168), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n706), .B2(G21), .ZN(new_n708));
  INV_X1    g283(.A(G1966), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2072), .ZN(new_n711));
  OR2_X1    g286(.A1(G29), .A2(G33), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n624), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(new_n478), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n472), .A2(G139), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT99), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT98), .B(KEYINPUT25), .Z(new_n719));
  NAND3_X1  g294(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n716), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n712), .B1(new_n723), .B2(new_n695), .ZN(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n695), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n695), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT29), .Z(new_n728));
  OAI221_X1 g303(.A(new_n710), .B1(new_n711), .B2(new_n724), .C1(new_n725), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n695), .A2(G32), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT26), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n473), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n732), .B(new_n734), .C1(G129), .C2(new_n479), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(new_n695), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT27), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G1996), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n724), .A2(new_n711), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n737), .A2(G1996), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n729), .A2(new_n738), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G171), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT103), .B(G1961), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n695), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n695), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2078), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n695), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n472), .A2(G140), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT96), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n479), .B2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT97), .B(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n743), .A2(new_n744), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n745), .A2(new_n748), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n708), .A2(new_n709), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT101), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n728), .A2(new_n725), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT104), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n741), .A2(new_n762), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT89), .B(G16), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n543), .B2(new_n769), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT95), .B(G1341), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n771), .B(new_n772), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n706), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n611), .B2(new_n706), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1348), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n768), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n580), .B2(new_n706), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n767), .A2(new_n773), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n595), .A2(new_n706), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G6), .B2(new_n706), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n706), .A2(G23), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G288), .B2(G16), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n783), .A2(new_n784), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n768), .A2(G22), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n768), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1971), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n783), .B2(new_n784), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n790), .A2(KEYINPUT34), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT34), .B1(new_n790), .B2(new_n795), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n768), .B1(G290), .B2(KEYINPUT91), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT91), .B2(G290), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n768), .A2(G24), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT90), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT92), .B(G1986), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n695), .A2(G25), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n472), .A2(G131), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n479), .A2(G119), .ZN(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n805), .B1(new_n811), .B2(new_n695), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n796), .A2(new_n797), .A3(new_n804), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n781), .A2(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n512), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n516), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n512), .A2(G93), .A3(new_n497), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n499), .A2(G55), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT107), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT106), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n611), .A2(G559), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n542), .A2(new_n825), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n821), .A2(new_n824), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(new_n536), .C1(new_n541), .C2(new_n540), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n839), .A2(KEYINPUT39), .A3(new_n840), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n829), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n840), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n833), .A2(new_n838), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  AND4_X1   g424(.A1(new_n829), .A2(new_n848), .A3(new_n849), .A4(new_n844), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n828), .B1(new_n845), .B2(new_n850), .ZN(G145));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n479), .A2(G126), .ZN(new_n853));
  INV_X1    g428(.A(new_n493), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT108), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT108), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n494), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n490), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n757), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n723), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(new_n735), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n479), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n478), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G142), .B2(new_n472), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n626), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n810), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n862), .A2(new_n869), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n475), .B(new_n636), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n483), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n873), .A2(new_n870), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n852), .B1(new_n877), .B2(new_n878), .C1(new_n876), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g456(.A(new_n619), .B(new_n837), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n580), .A2(new_n610), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n567), .A2(new_n579), .A3(new_n609), .A4(new_n606), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  AND4_X1   g462(.A1(new_n567), .A2(new_n579), .A3(new_n609), .A4(new_n606), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n567), .A2(new_n579), .B1(new_n606), .B2(new_n609), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(KEYINPUT41), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT42), .Z(new_n895));
  OAI211_X1 g470(.A(new_n586), .B(new_n588), .C1(new_n591), .C2(new_n594), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n598), .B2(new_n599), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n598), .A2(new_n599), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(G166), .A2(KEYINPUT111), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(G166), .A2(KEYINPUT111), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n899), .B(new_n900), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n595), .A2(G288), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n906));
  NAND2_X1  g481(.A1(G303), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n900), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n907), .B(new_n901), .C1(new_n908), .C2(new_n898), .ZN(new_n909));
  AND4_X1   g484(.A1(new_n896), .A2(new_n904), .A3(new_n905), .A4(new_n909), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n909), .A2(new_n904), .B1(new_n905), .B2(new_n896), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n895), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n895), .A2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n825), .A2(new_n601), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n834), .A2(G301), .A3(new_n836), .ZN(new_n920));
  AOI21_X1  g495(.A(G301), .B1(new_n834), .B2(new_n836), .ZN(new_n921));
  OAI21_X1  g496(.A(G286), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n542), .A2(new_n825), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n537), .A2(new_n539), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT74), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n537), .A2(KEYINPUT74), .A3(new_n539), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n835), .B1(new_n928), .B2(new_n536), .ZN(new_n929));
  OAI21_X1  g504(.A(G171), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n834), .A2(new_n836), .A3(G301), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(G168), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n892), .A2(new_n922), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n892), .A2(new_n922), .A3(new_n932), .A4(KEYINPUT112), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n920), .A2(new_n921), .A3(G286), .ZN(new_n937));
  AOI21_X1  g512(.A(G168), .B1(new_n930), .B2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n885), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n935), .A2(new_n912), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n852), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n912), .B1(new_n942), .B2(KEYINPUT113), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n935), .A2(new_n944), .A3(new_n936), .A4(new_n939), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n919), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n937), .A2(new_n938), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n939), .A2(KEYINPUT114), .B1(new_n949), .B2(new_n892), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n922), .A2(new_n932), .B1(new_n883), .B2(new_n884), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n912), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT115), .B1(new_n954), .B2(new_n941), .ZN(new_n955));
  INV_X1    g530(.A(new_n912), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n933), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n939), .A2(KEYINPUT114), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n852), .A4(new_n940), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n948), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(KEYINPUT113), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n956), .A3(new_n945), .ZN(new_n965));
  INV_X1    g540(.A(new_n941), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n947), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n954), .A2(new_n941), .A3(KEYINPUT43), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n919), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n963), .A2(KEYINPUT116), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n859), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(G160), .A2(G40), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  INV_X1    g560(.A(G2067), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n757), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n979), .B1(new_n987), .B2(new_n735), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n983), .B2(new_n982), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n735), .B(G1996), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(new_n987), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n811), .A2(new_n813), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n811), .A2(new_n813), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n979), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n979), .A2(G1986), .A3(G290), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(KEYINPUT48), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(KEYINPUT48), .B2(new_n998), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n994), .B(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G2067), .B2(new_n757), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n980), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n991), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n859), .A2(new_n975), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n977), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(G288), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  INV_X1    g587(.A(G288), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(G1976), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(KEYINPUT52), .B2(new_n1011), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n495), .A2(new_n975), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n859), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n978), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(G1971), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(new_n978), .C1(KEYINPUT50), .C2(new_n1006), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(G2090), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1008), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G166), .A2(new_n1008), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT55), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1009), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n591), .A2(G1981), .A3(new_n594), .ZN(new_n1031));
  INV_X1    g606(.A(new_n590), .ZN(new_n1032));
  OAI21_X1  g607(.A(G1981), .B1(new_n1032), .B2(new_n594), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(KEYINPUT117), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1016), .B(new_n1029), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n977), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1022), .B1(G2090), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1028), .B1(new_n1045), .B2(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n976), .B2(new_n977), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  AOI22_X1  g623(.A1(KEYINPUT108), .A2(new_n855), .B1(new_n487), .B2(new_n489), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n858), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1048), .B(new_n978), .C1(new_n1050), .C2(KEYINPUT45), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n709), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1024), .A2(G2084), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1008), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G168), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1040), .A2(new_n1046), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT63), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1059), .A2(new_n1057), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1058), .A2(KEYINPUT63), .B1(new_n1040), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1016), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1062), .A2(new_n1029), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1031), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1009), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1956), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT56), .B(G2072), .Z(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT119), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1021), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT57), .B1(new_n553), .B2(new_n566), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n578), .A2(new_n1075), .A3(new_n550), .A4(new_n568), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1070), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1070), .A2(KEYINPUT120), .A3(new_n1073), .A4(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1073), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1077), .B1(new_n1084), .B2(new_n1069), .ZN(new_n1085));
  INV_X1    g660(.A(G1348), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1024), .A2(new_n1086), .B1(new_n986), .B2(new_n1007), .ZN(new_n1087));
  INV_X1    g662(.A(new_n611), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1019), .A2(new_n981), .A3(new_n1020), .A4(new_n978), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1007), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n543), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT59), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1085), .A2(new_n1079), .A3(KEYINPUT61), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  OR3_X1    g673(.A1(new_n1087), .A2(new_n1088), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1088), .A2(new_n1098), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1087), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1090), .B1(new_n1091), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G286), .A2(G8), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT121), .Z(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT51), .B1(new_n1056), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT122), .B(KEYINPUT51), .C1(new_n1056), .C2(new_n1106), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1105), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1056), .A2(KEYINPUT51), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G2078), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n1021), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1961), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1024), .ZN(new_n1120));
  XOR2_X1   g695(.A(G301), .B(KEYINPUT54), .Z(new_n1121));
  OR3_X1    g696(.A1(new_n976), .A2(KEYINPUT124), .A3(new_n977), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n976), .B2(new_n977), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n1117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1120), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1053), .A2(G2078), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT53), .B1(new_n1127), .B2(KEYINPUT123), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1120), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1121), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1104), .A2(new_n1116), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT125), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1113), .A2(new_n1135), .A3(new_n1115), .ZN(new_n1136));
  AOI21_X1  g711(.A(G301), .B1(KEYINPUT125), .B2(new_n1134), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1130), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1133), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1068), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(G290), .B(G1986), .Z(new_n1144));
  AOI21_X1  g719(.A(new_n979), .B1(new_n996), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1005), .B1(new_n1143), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g721(.A1(new_n967), .A2(new_n968), .ZN(new_n1148));
  NOR4_X1   g722(.A1(G229), .A2(G401), .A3(new_n460), .A4(G227), .ZN(new_n1149));
  NAND3_X1  g723(.A1(new_n880), .A2(new_n1148), .A3(new_n1149), .ZN(G225));
  INV_X1    g724(.A(G225), .ZN(G308));
endmodule


