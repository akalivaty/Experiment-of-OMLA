//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(new_n463), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n474), .A2(KEYINPUT64), .A3(G124), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n477), .A2(new_n479), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT65), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n473), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n460), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n490));
  NOR2_X1   g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n473), .B2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(new_n494), .B2(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(new_n463), .A3(G126), .A4(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n487), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n500), .A2(KEYINPUT6), .A3(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT6), .B1(new_n500), .B2(G651), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n501), .A2(new_n502), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n508), .A2(new_n510), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G62), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n506), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NOR2_X1   g093(.A1(new_n507), .A2(new_n505), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n512), .A2(G90), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(G52), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n511), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n519), .A2(G43), .B1(G651), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n512), .A2(G81), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n503), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n548), .A2(KEYINPUT9), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n548), .B2(new_n549), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(new_n551), .B1(G91), .B2(new_n512), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n529), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT69), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  NAND2_X1  g132(.A1(new_n519), .A2(G49), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n512), .A2(G87), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  AOI22_X1  g136(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n529), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n512), .A2(KEYINPUT71), .A3(G86), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n512), .A2(G86), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(new_n568), .B1(G48), .B2(new_n519), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n565), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(G305));
  NAND2_X1  g146(.A1(new_n512), .A2(G85), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n519), .A2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n529), .C2(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G171), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n505), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(G54), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n529), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n582), .A2(KEYINPUT74), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT74), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n512), .A2(G92), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT10), .Z(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT72), .B1(new_n590), .B2(new_n576), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n579), .B1(new_n591), .B2(new_n577), .ZN(G284));
  OAI21_X1  g167(.A(new_n579), .B1(new_n591), .B2(new_n577), .ZN(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  XOR2_X1   g169(.A(G299), .B(KEYINPUT75), .Z(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  AND2_X1   g172(.A1(new_n587), .A2(new_n589), .ZN(new_n598));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n478), .A2(G2104), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  INV_X1    g185(.A(G123), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n475), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n478), .A2(G135), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT78), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT78), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n615), .B(new_n616), .C1(G111), .C2(new_n473), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n474), .A2(KEYINPUT77), .A3(G123), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n612), .A2(new_n613), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n609), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2438), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2443), .B(G2446), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n634), .A2(G14), .ZN(G401));
  XNOR2_X1  g210(.A(G2072), .B(G2078), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2084), .B(G2090), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n638), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(new_n636), .B2(new_n639), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT80), .Z(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n640), .B2(new_n638), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n639), .A3(new_n636), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT79), .B(KEYINPUT18), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n620), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(KEYINPUT20), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n662), .A3(new_n659), .ZN(new_n669));
  NAND4_X1  g244(.A1(new_n664), .A2(new_n665), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT86), .B(G1986), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G29), .B2(G33), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n678), .A2(G29), .A3(G33), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n478), .A2(G139), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT94), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n473), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT25), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n679), .B(new_n680), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2072), .ZN(new_n690));
  INV_X1    g265(.A(G2084), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT95), .ZN(new_n692));
  NOR2_X1   g267(.A1(KEYINPUT24), .A2(G34), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(KEYINPUT24), .A2(G34), .ZN(new_n695));
  AOI21_X1  g270(.A(G29), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g271(.A1(G160), .A2(G29), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n692), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G32), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n468), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G2105), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n474), .A2(G129), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT96), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT96), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  AND3_X1   g282(.A1(new_n705), .A2(KEYINPUT97), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(KEYINPUT97), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n699), .B1(new_n711), .B2(new_n688), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT27), .B(G1996), .Z(new_n713));
  OAI221_X1 g288(.A(new_n690), .B1(new_n691), .B2(new_n698), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT98), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n688), .A2(G35), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G162), .B2(new_n688), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT100), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT29), .B(G2090), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(KEYINPUT30), .A2(G28), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT30), .A2(G28), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n721), .A2(new_n722), .A3(G29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n619), .B2(G29), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n712), .B2(new_n713), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n688), .A2(G26), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n727));
  INV_X1    g302(.A(G104), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n473), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n474), .A2(G128), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n478), .A2(G140), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n726), .B1(new_n734), .B2(new_n688), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n726), .B(new_n735), .S(KEYINPUT28), .Z(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G19), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n541), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  INV_X1    g318(.A(G1341), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n725), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n691), .B2(new_n698), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n740), .A2(KEYINPUT23), .A3(G20), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT23), .B1(new_n740), .B2(G20), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n748), .B(new_n749), .C1(G299), .C2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1956), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n688), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n688), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n755), .C1(new_n744), .C2(new_n743), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n715), .A2(new_n720), .A3(new_n747), .A4(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G16), .A2(G21), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G168), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT99), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n765));
  MUX2_X1   g340(.A(G6), .B(G305), .S(G16), .Z(new_n766));
  XOR2_X1   g341(.A(KEYINPUT32), .B(G1981), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT89), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n740), .A2(G22), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G166), .B2(new_n740), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1971), .Z(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G23), .ZN(new_n773));
  INV_X1    g348(.A(G288), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT33), .B(G1976), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n769), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT34), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT34), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n780), .A2(new_n784), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n688), .A2(G25), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n788));
  INV_X1    g363(.A(G95), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n473), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT87), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G131), .B2(new_n478), .ZN(new_n792));
  INV_X1    g367(.A(G119), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n475), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT88), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n798), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n740), .A2(G24), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G290), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1986), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n799), .A2(new_n800), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n765), .B1(new_n786), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g383(.A(KEYINPUT36), .B(new_n806), .C1(new_n783), .C2(new_n785), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n759), .B(new_n764), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n740), .A2(G5), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G171), .B2(new_n740), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1961), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n740), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n598), .B2(new_n740), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n810), .A2(new_n813), .A3(new_n818), .ZN(G311));
  INV_X1    g394(.A(new_n808), .ZN(new_n820));
  INV_X1    g395(.A(new_n809), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n758), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n813), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n817), .A4(new_n764), .ZN(G150));
  NAND2_X1  g399(.A1(new_n512), .A2(G93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n519), .A2(G55), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n825), .B(new_n826), .C1(new_n529), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n541), .B(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n599), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT101), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  INV_X1    g413(.A(G37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n705), .A2(new_n707), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n490), .B1(new_n489), .B2(new_n492), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n494), .A2(KEYINPUT66), .A3(new_n491), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n497), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n496), .A2(new_n846), .A3(new_n497), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n841), .B1(new_n848), .B2(new_n487), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT4), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n486), .B(new_n850), .ZN(new_n851));
  AOI211_X1 g426(.A(KEYINPUT104), .B(new_n851), .C1(new_n845), .C2(new_n847), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n733), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n496), .A2(new_n846), .A3(new_n497), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n846), .B1(new_n496), .B2(new_n497), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n487), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n848), .A2(new_n841), .A3(new_n487), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n734), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n854), .B1(new_n853), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n840), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n849), .A2(new_n852), .A3(new_n733), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n734), .B1(new_n858), .B2(new_n859), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT105), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n840), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n687), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n711), .A2(new_n853), .A3(new_n860), .ZN(new_n871));
  INV_X1    g446(.A(new_n687), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n710), .B1(new_n864), .B2(new_n865), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n474), .A2(G130), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n478), .A2(G142), .ZN(new_n877));
  NOR2_X1   g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n607), .B(new_n880), .Z(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n794), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n470), .B(KEYINPUT102), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n484), .B(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n619), .Z(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n870), .A2(new_n874), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n870), .B2(new_n874), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n890), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n839), .B(new_n889), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  INV_X1    g474(.A(new_n888), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n870), .B2(new_n874), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n901), .A3(new_n892), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n875), .A2(new_n892), .A3(new_n882), .ZN(new_n903));
  INV_X1    g478(.A(new_n886), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(KEYINPUT108), .A3(new_n839), .A4(new_n889), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT40), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n898), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(G395));
  NAND2_X1  g489(.A1(new_n828), .A2(new_n576), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G288), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(G305), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(G305), .ZN(new_n918));
  XOR2_X1   g493(.A(G290), .B(KEYINPUT109), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(KEYINPUT110), .B2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n598), .B(G299), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n590), .B(G299), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT41), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n601), .B(new_n829), .ZN(new_n930));
  MUX2_X1   g505(.A(new_n927), .B(new_n929), .S(new_n930), .Z(new_n931));
  XNOR2_X1  g506(.A(new_n926), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n915), .B1(new_n932), .B2(new_n576), .ZN(G295));
  OAI21_X1  g508(.A(new_n915), .B1(new_n932), .B2(new_n576), .ZN(G331));
  XNOR2_X1  g509(.A(new_n829), .B(G286), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(G171), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n928), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n927), .A2(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n940), .A3(new_n936), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n941), .B2(KEYINPUT112), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n929), .A2(new_n943), .A3(new_n936), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n923), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n928), .B2(new_n936), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n921), .A2(KEYINPUT113), .A3(new_n922), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT113), .B1(new_n921), .B2(new_n922), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n839), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n839), .ZN(new_n953));
  INV_X1    g528(.A(new_n949), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n944), .B2(new_n942), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(KEYINPUT44), .B(new_n952), .C1(new_n956), .C2(KEYINPUT43), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n953), .B2(new_n955), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n945), .A2(new_n959), .A3(new_n839), .A4(new_n950), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(G397));
  NAND2_X1  g539(.A1(new_n858), .A2(new_n859), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT114), .B(G1384), .Z(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G160), .A2(G40), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT48), .Z(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n867), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n733), .B(G2067), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n976), .B(new_n977), .C1(new_n711), .C2(new_n975), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n794), .B(new_n798), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n974), .B1(new_n971), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n971), .B1(new_n840), .B2(new_n977), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(KEYINPUT46), .A3(new_n975), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n970), .B2(G1996), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  NOR2_X1   g562(.A1(new_n794), .A2(new_n797), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n978), .A2(new_n988), .B1(new_n737), .B2(new_n734), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n970), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n981), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(G305), .A2(G1981), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n519), .A2(G48), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n563), .A2(new_n567), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G1981), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(KEYINPUT118), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(KEYINPUT118), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n992), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n851), .B1(new_n845), .B2(new_n847), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1001), .A2(KEYINPUT116), .A3(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n857), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n969), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n992), .A2(new_n996), .A3(KEYINPUT49), .A4(new_n997), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1000), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n774), .A2(G1976), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  OR3_X1    g589(.A1(new_n1013), .A2(KEYINPUT117), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT117), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1014), .C1(G1976), .C2(new_n774), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT115), .B(G1971), .Z(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n966), .C1(new_n849), .C2(new_n852), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1021), .A2(G40), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n498), .A2(new_n1004), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n470), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1020), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1023), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n969), .B1(new_n1029), .B2(new_n1027), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2090), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n1008), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT55), .Z(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1011), .A2(G1976), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n992), .B1(new_n1040), .B2(G288), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1019), .A2(new_n1039), .B1(new_n1041), .B2(new_n1009), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1017), .A2(new_n1038), .A3(KEYINPUT63), .A4(new_n1018), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT116), .B1(new_n1001), .B2(G1384), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n857), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT50), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1046), .A2(G2084), .A3(new_n1030), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1024), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT45), .B(new_n1004), .C1(new_n851), .C2(new_n844), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n498), .A2(KEYINPUT120), .A3(KEYINPUT45), .A4(new_n1004), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n968), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1966), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n1043), .A2(G286), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1042), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n763), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1028), .A2(new_n1031), .A3(new_n691), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1008), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G286), .A2(G8), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT123), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1060), .B(new_n1061), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1067), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1071));
  NAND2_X1  g646(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1055), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT125), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1022), .A2(new_n754), .A3(new_n1025), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(new_n1032), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n754), .A2(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1062), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1075), .A2(new_n1086), .A3(new_n1077), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1079), .A2(G171), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1021), .A2(G40), .A3(new_n975), .A4(new_n1025), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1006), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT122), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1093), .A2(KEYINPUT59), .A3(new_n541), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n816), .B1(new_n1046), .B2(new_n1030), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n737), .B(new_n969), .C1(new_n1002), .C2(new_n1005), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1097), .A2(new_n590), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n590), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n598), .A2(new_n1097), .A3(new_n1102), .A4(new_n1098), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1096), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1093), .A2(new_n541), .A3(new_n1095), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G299), .B(KEYINPUT57), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1021), .A2(G40), .A3(new_n1025), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT50), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n968), .B1(new_n1029), .B2(new_n1027), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1107), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G299), .B(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(new_n1109), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1105), .A2(new_n1106), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1114), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1104), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1115), .B2(new_n1109), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1124), .B2(new_n1100), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G171), .B(KEYINPUT54), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n469), .A2(G2105), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n967), .A2(new_n1129), .A3(new_n1084), .ZN(new_n1130));
  INV_X1    g705(.A(new_n466), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n473), .B1(new_n1131), .B2(KEYINPUT126), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(KEYINPUT126), .B2(new_n1131), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1022), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1083), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1128), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1085), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1127), .A2(new_n1078), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(G168), .B(new_n1065), .C1(new_n1043), .C2(new_n1056), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1088), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1019), .A2(new_n1038), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G2090), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1026), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1008), .B1(new_n1144), .B2(KEYINPUT119), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1037), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1059), .B1(new_n1140), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(G290), .A2(G1986), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n980), .A2(new_n972), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n970), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n991), .B1(new_n1149), .B2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g728(.A(G319), .ZN(new_n1155));
  OR2_X1    g729(.A1(G227), .A2(new_n1155), .ZN(new_n1156));
  OR2_X1    g730(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1157));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1158));
  NOR3_X1   g732(.A1(new_n1158), .A2(G229), .A3(G401), .ZN(new_n1159));
  AND4_X1   g733(.A1(new_n910), .A2(new_n961), .A3(new_n1157), .A4(new_n1159), .ZN(G308));
  NAND4_X1  g734(.A1(new_n910), .A2(new_n961), .A3(new_n1157), .A4(new_n1159), .ZN(G225));
endmodule


