

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788;

  AND2_X1 U381 ( .A1(n767), .A2(n391), .ZN(n708) );
  AND2_X1 U382 ( .A1(n689), .A2(n574), .ZN(n403) );
  NOR2_X1 U383 ( .A1(n641), .A2(n765), .ZN(n366) );
  BUF_X1 U384 ( .A(n711), .Z(n362) );
  INV_X1 U385 ( .A(n617), .ZN(n360) );
  NAND2_X1 U386 ( .A1(n364), .A2(n363), .ZN(n632) );
  INV_X1 U387 ( .A(n729), .ZN(n363) );
  INV_X1 U388 ( .A(n627), .ZN(n364) );
  XNOR2_X1 U389 ( .A(n542), .B(KEYINPUT0), .ZN(n594) );
  NAND2_X1 U390 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U391 ( .A(n525), .B(KEYINPUT107), .ZN(n727) );
  OR2_X1 U392 ( .A1(n564), .A2(n714), .ZN(n566) );
  NAND2_X1 U393 ( .A1(n400), .A2(n397), .ZN(n608) );
  NAND2_X1 U394 ( .A1(n405), .A2(n408), .ZN(n622) );
  XNOR2_X1 U395 ( .A(n484), .B(n772), .ZN(n671) );
  XNOR2_X1 U396 ( .A(n479), .B(n376), .ZN(n470) );
  XNOR2_X1 U397 ( .A(n365), .B(KEYINPUT71), .ZN(n499) );
  INV_X1 U398 ( .A(G131), .ZN(n365) );
  XNOR2_X2 U399 ( .A(n361), .B(n360), .ZN(n646) );
  NAND2_X1 U400 ( .A1(n630), .A2(n615), .ZN(n361) );
  NAND2_X2 U401 ( .A1(n416), .A2(n414), .ZN(n573) );
  OR2_X2 U402 ( .A1(n611), .A2(n551), .ZN(n462) );
  NAND2_X1 U403 ( .A1(n643), .A2(n366), .ZN(n644) );
  NAND2_X2 U404 ( .A1(n563), .A2(n562), .ZN(n587) );
  XNOR2_X1 U405 ( .A(G119), .B(G128), .ZN(n440) );
  AND2_X2 U406 ( .A1(n614), .A2(n613), .ZN(n630) );
  AND2_X2 U407 ( .A1(n571), .A2(n572), .ZN(n525) );
  INV_X2 U408 ( .A(G953), .ZN(n782) );
  INV_X1 U409 ( .A(n372), .ZN(n688) );
  AND2_X1 U410 ( .A1(n419), .A2(n417), .ZN(n416) );
  XNOR2_X1 U411 ( .A(n470), .B(n435), .ZN(n666) );
  INV_X1 U412 ( .A(KEYINPUT40), .ZN(n374) );
  XNOR2_X1 U413 ( .A(G125), .B(KEYINPUT10), .ZN(n413) );
  XNOR2_X1 U414 ( .A(n375), .B(n374), .ZN(n687) );
  AND2_X1 U415 ( .A1(n631), .A2(n757), .ZN(n640) );
  OR2_X1 U416 ( .A1(n367), .A2(n627), .ZN(n631) );
  NAND2_X2 U417 ( .A1(n388), .A2(n384), .ZN(n546) );
  AND2_X1 U418 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U419 ( .A(n470), .B(n469), .ZN(n700) );
  XNOR2_X1 U420 ( .A(n413), .B(G146), .ZN(n495) );
  OR2_X1 U421 ( .A1(n729), .A2(KEYINPUT47), .ZN(n367) );
  NAND2_X1 U422 ( .A1(n622), .A2(n490), .ZN(n370) );
  NAND2_X1 U423 ( .A1(n368), .A2(n369), .ZN(n371) );
  NAND2_X1 U424 ( .A1(n370), .A2(n371), .ZN(n541) );
  INV_X1 U425 ( .A(n622), .ZN(n368) );
  INV_X1 U426 ( .A(n490), .ZN(n369) );
  XOR2_X1 U427 ( .A(n462), .B(KEYINPUT28), .Z(n425) );
  XNOR2_X1 U428 ( .A(n373), .B(KEYINPUT32), .ZN(n372) );
  NOR2_X1 U429 ( .A1(n585), .A2(n584), .ZN(n373) );
  AND2_X1 U430 ( .A1(n402), .A2(n401), .ZN(n400) );
  NOR2_X2 U431 ( .A1(n646), .A2(n760), .ZN(n375) );
  NOR2_X2 U432 ( .A1(n705), .A2(n393), .ZN(n392) );
  AND2_X2 U433 ( .A1(n607), .A2(n711), .ZN(n595) );
  XNOR2_X1 U434 ( .A(n507), .B(G475), .ZN(n572) );
  INV_X1 U435 ( .A(KEYINPUT2), .ZN(n393) );
  NAND2_X1 U436 ( .A1(n486), .A2(n651), .ZN(n411) );
  NAND2_X1 U437 ( .A1(n410), .A2(n649), .ZN(n409) );
  INV_X1 U438 ( .A(n486), .ZN(n410) );
  OR2_X1 U439 ( .A1(n666), .A2(n385), .ZN(n384) );
  NAND2_X1 U440 ( .A1(n387), .A2(n386), .ZN(n385) );
  OR2_X1 U441 ( .A1(n700), .A2(n398), .ZN(n397) );
  NAND2_X1 U442 ( .A1(n399), .A2(n386), .ZN(n398) );
  XOR2_X1 U443 ( .A(G137), .B(G140), .Z(n463) );
  XNOR2_X1 U444 ( .A(n644), .B(n423), .ZN(n648) );
  NOR2_X1 U445 ( .A1(n418), .A2(n628), .ZN(n417) );
  NOR2_X1 U446 ( .A1(n569), .A2(n570), .ZN(n418) );
  XNOR2_X1 U447 ( .A(n499), .B(n428), .ZN(n777) );
  XNOR2_X1 U448 ( .A(n421), .B(n420), .ZN(n679) );
  XNOR2_X1 U449 ( .A(n445), .B(n439), .ZN(n420) );
  XNOR2_X1 U450 ( .A(n443), .B(n778), .ZN(n421) );
  XNOR2_X1 U451 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U452 ( .A(n502), .B(n422), .ZN(n503) );
  AND2_X1 U453 ( .A1(n406), .A2(n381), .ZN(n405) );
  INV_X1 U454 ( .A(n724), .ZN(n407) );
  BUF_X1 U455 ( .A(n564), .Z(n713) );
  NAND2_X1 U456 ( .A1(n415), .A2(KEYINPUT34), .ZN(n414) );
  XOR2_X1 U457 ( .A(n777), .B(G146), .Z(n376) );
  OR2_X1 U458 ( .A1(n689), .A2(n576), .ZN(n377) );
  OR2_X1 U459 ( .A1(n586), .A2(n372), .ZN(n378) );
  AND2_X1 U460 ( .A1(n569), .A2(n570), .ZN(n379) );
  AND2_X1 U461 ( .A1(n604), .A2(n603), .ZN(n380) );
  AND2_X1 U462 ( .A1(n407), .A2(n411), .ZN(n381) );
  INV_X1 U463 ( .A(G902), .ZN(n386) );
  XOR2_X1 U464 ( .A(KEYINPUT90), .B(KEYINPUT35), .Z(n382) );
  XOR2_X1 U465 ( .A(n605), .B(KEYINPUT64), .Z(n383) );
  NAND2_X1 U466 ( .A1(n666), .A2(n436), .ZN(n390) );
  XNOR2_X2 U467 ( .A(n546), .B(KEYINPUT109), .ZN(n611) );
  INV_X1 U468 ( .A(n436), .ZN(n387) );
  NAND2_X1 U469 ( .A1(n436), .A2(G902), .ZN(n389) );
  XNOR2_X1 U470 ( .A(n392), .B(n656), .ZN(n391) );
  XNOR2_X2 U471 ( .A(n394), .B(n383), .ZN(n767) );
  NAND2_X1 U472 ( .A1(n395), .A2(n380), .ZN(n394) );
  NAND2_X1 U473 ( .A1(n396), .A2(n377), .ZN(n395) );
  NAND2_X1 U474 ( .A1(n403), .A2(n378), .ZN(n396) );
  NAND2_X1 U475 ( .A1(n700), .A2(n472), .ZN(n402) );
  XNOR2_X2 U476 ( .A(n608), .B(KEYINPUT1), .ZN(n711) );
  INV_X1 U477 ( .A(n472), .ZN(n399) );
  NAND2_X1 U478 ( .A1(n472), .A2(G902), .ZN(n401) );
  NAND2_X1 U479 ( .A1(n404), .A2(n408), .ZN(n526) );
  OR2_X1 U480 ( .A1(n671), .A2(n409), .ZN(n408) );
  AND2_X1 U481 ( .A1(n406), .A2(n411), .ZN(n404) );
  NAND2_X1 U482 ( .A1(n671), .A2(n486), .ZN(n406) );
  XNOR2_X2 U483 ( .A(n412), .B(G143), .ZN(n516) );
  XNOR2_X2 U484 ( .A(G128), .B(KEYINPUT66), .ZN(n412) );
  INV_X1 U485 ( .A(n733), .ZN(n415) );
  NAND2_X1 U486 ( .A1(n733), .A2(n379), .ZN(n419) );
  XNOR2_X2 U487 ( .A(n568), .B(KEYINPUT33), .ZN(n733) );
  BUF_X1 U488 ( .A(n692), .Z(n697) );
  AND2_X2 U489 ( .A1(n697), .A2(G478), .ZN(n693) );
  XNOR2_X1 U490 ( .A(n504), .B(n503), .ZN(n658) );
  XNOR2_X1 U491 ( .A(n479), .B(n478), .ZN(n484) );
  XOR2_X1 U492 ( .A(n501), .B(n500), .Z(n422) );
  XOR2_X1 U493 ( .A(KEYINPUT72), .B(KEYINPUT48), .Z(n423) );
  AND2_X1 U494 ( .A1(n647), .A2(n686), .ZN(n424) );
  INV_X1 U495 ( .A(KEYINPUT105), .ZN(n510) );
  INV_X1 U496 ( .A(KEYINPUT89), .ZN(n656) );
  INV_X1 U497 ( .A(KEYINPUT34), .ZN(n570) );
  XNOR2_X1 U498 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U499 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X2 U500 ( .A(n516), .B(n426), .ZN(n781) );
  XNOR2_X2 U501 ( .A(n781), .B(G101), .ZN(n479) );
  INV_X1 U502 ( .A(G134), .ZN(n428) );
  NOR2_X1 U503 ( .A1(G953), .A2(G237), .ZN(n494) );
  NAND2_X1 U504 ( .A1(n494), .A2(G210), .ZN(n429) );
  XNOR2_X1 U505 ( .A(n429), .B(G137), .ZN(n431) );
  XNOR2_X1 U506 ( .A(KEYINPUT79), .B(KEYINPUT5), .ZN(n430) );
  XNOR2_X1 U507 ( .A(n431), .B(n430), .ZN(n434) );
  XNOR2_X1 U508 ( .A(G113), .B(G116), .ZN(n433) );
  XNOR2_X1 U509 ( .A(KEYINPUT3), .B(G119), .ZN(n432) );
  XNOR2_X1 U510 ( .A(n433), .B(n432), .ZN(n482) );
  XNOR2_X1 U511 ( .A(n434), .B(n482), .ZN(n435) );
  XNOR2_X1 U512 ( .A(KEYINPUT98), .B(G472), .ZN(n436) );
  XOR2_X1 U513 ( .A(n495), .B(n463), .Z(n778) );
  XOR2_X1 U514 ( .A(KEYINPUT95), .B(KEYINPUT86), .Z(n438) );
  XNOR2_X1 U515 ( .A(G110), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U516 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U517 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n441) );
  XNOR2_X1 U518 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U519 ( .A(n442), .B(KEYINPUT23), .Z(n443) );
  NAND2_X1 U520 ( .A1(G234), .A2(n782), .ZN(n444) );
  XOR2_X1 U521 ( .A(KEYINPUT8), .B(n444), .Z(n515) );
  AND2_X1 U522 ( .A1(n515), .A2(G221), .ZN(n445) );
  NAND2_X1 U523 ( .A1(n679), .A2(n386), .ZN(n449) );
  XNOR2_X1 U524 ( .A(KEYINPUT15), .B(G902), .ZN(n649) );
  NAND2_X1 U525 ( .A1(n649), .A2(G234), .ZN(n446) );
  XNOR2_X1 U526 ( .A(n446), .B(KEYINPUT20), .ZN(n450) );
  NAND2_X1 U527 ( .A1(n450), .A2(G217), .ZN(n447) );
  XNOR2_X1 U528 ( .A(n447), .B(KEYINPUT25), .ZN(n448) );
  XNOR2_X1 U529 ( .A(n449), .B(n448), .ZN(n564) );
  XOR2_X1 U530 ( .A(KEYINPUT21), .B(KEYINPUT97), .Z(n452) );
  NAND2_X1 U531 ( .A1(n450), .A2(G221), .ZN(n451) );
  XNOR2_X1 U532 ( .A(n452), .B(n451), .ZN(n714) );
  NAND2_X1 U533 ( .A1(G953), .A2(G902), .ZN(n534) );
  NOR2_X1 U534 ( .A1(G900), .A2(n534), .ZN(n454) );
  NAND2_X1 U535 ( .A1(G237), .A2(G234), .ZN(n453) );
  XNOR2_X1 U536 ( .A(n453), .B(KEYINPUT14), .ZN(n738) );
  AND2_X1 U537 ( .A1(n454), .A2(n738), .ZN(n456) );
  INV_X1 U538 ( .A(KEYINPUT112), .ZN(n455) );
  XNOR2_X1 U539 ( .A(n456), .B(n455), .ZN(n459) );
  NAND2_X1 U540 ( .A1(n782), .A2(G952), .ZN(n538) );
  INV_X1 U541 ( .A(n538), .ZN(n457) );
  NAND2_X1 U542 ( .A1(n738), .A2(n457), .ZN(n458) );
  NAND2_X1 U543 ( .A1(n459), .A2(n458), .ZN(n606) );
  INV_X1 U544 ( .A(n606), .ZN(n460) );
  NOR2_X1 U545 ( .A1(n714), .A2(n460), .ZN(n461) );
  NAND2_X1 U546 ( .A1(n564), .A2(n461), .ZN(n551) );
  XOR2_X1 U547 ( .A(n463), .B(KEYINPUT81), .Z(n468) );
  XNOR2_X1 U548 ( .A(G107), .B(G104), .ZN(n465) );
  XNOR2_X1 U549 ( .A(KEYINPUT93), .B(G110), .ZN(n464) );
  XNOR2_X1 U550 ( .A(n465), .B(n464), .ZN(n481) );
  NAND2_X1 U551 ( .A1(G227), .A2(n782), .ZN(n466) );
  XNOR2_X1 U552 ( .A(n481), .B(n466), .ZN(n467) );
  XNOR2_X1 U553 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U554 ( .A(KEYINPUT73), .ZN(n471) );
  XNOR2_X1 U555 ( .A(n471), .B(G469), .ZN(n472) );
  NAND2_X1 U556 ( .A1(n425), .A2(n608), .ZN(n529) );
  INV_X1 U557 ( .A(n529), .ZN(n491) );
  NAND2_X1 U558 ( .A1(n782), .A2(G224), .ZN(n473) );
  XNOR2_X1 U559 ( .A(n473), .B(KEYINPUT82), .ZN(n475) );
  XNOR2_X1 U560 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n474) );
  XNOR2_X1 U561 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U562 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U563 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U564 ( .A(KEYINPUT16), .B(G122), .ZN(n480) );
  XNOR2_X1 U565 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U566 ( .A(n483), .B(n482), .ZN(n772) );
  INV_X1 U567 ( .A(n649), .ZN(n651) );
  OR2_X1 U568 ( .A1(G237), .A2(G902), .ZN(n485) );
  XNOR2_X1 U569 ( .A(KEYINPUT78), .B(n485), .ZN(n487) );
  NAND2_X1 U570 ( .A1(n487), .A2(G210), .ZN(n486) );
  AND2_X1 U571 ( .A1(n487), .A2(G214), .ZN(n724) );
  XNOR2_X1 U572 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n489) );
  INV_X1 U573 ( .A(KEYINPUT69), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U575 ( .A1(n491), .A2(n541), .ZN(n627) );
  XOR2_X1 U576 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n493) );
  XNOR2_X1 U577 ( .A(G113), .B(KEYINPUT12), .ZN(n492) );
  XNOR2_X1 U578 ( .A(n493), .B(n492), .ZN(n498) );
  NAND2_X1 U579 ( .A1(G214), .A2(n494), .ZN(n496) );
  XNOR2_X1 U580 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U581 ( .A(n498), .B(n497), .Z(n504) );
  XNOR2_X1 U582 ( .A(n499), .B(KEYINPUT11), .ZN(n502) );
  XOR2_X1 U583 ( .A(G140), .B(G104), .Z(n501) );
  XNOR2_X1 U584 ( .A(G143), .B(G122), .ZN(n500) );
  NOR2_X1 U585 ( .A1(G902), .A2(n658), .ZN(n506) );
  XNOR2_X1 U586 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n505) );
  XNOR2_X1 U587 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U588 ( .A(n572), .B(KEYINPUT102), .ZN(n550) );
  XOR2_X1 U589 ( .A(G107), .B(KEYINPUT103), .Z(n509) );
  XNOR2_X1 U590 ( .A(G134), .B(KEYINPUT7), .ZN(n508) );
  XNOR2_X1 U591 ( .A(n509), .B(n508), .ZN(n513) );
  XNOR2_X1 U592 ( .A(G122), .B(KEYINPUT9), .ZN(n511) );
  XOR2_X1 U593 ( .A(n514), .B(KEYINPUT104), .Z(n520) );
  NAND2_X1 U594 ( .A1(n515), .A2(G217), .ZN(n518) );
  XNOR2_X1 U595 ( .A(n516), .B(G116), .ZN(n517) );
  XNOR2_X1 U596 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U597 ( .A(n520), .B(n519), .ZN(n694) );
  NAND2_X1 U598 ( .A1(n694), .A2(n386), .ZN(n522) );
  INV_X1 U599 ( .A(G478), .ZN(n521) );
  XNOR2_X1 U600 ( .A(n522), .B(n521), .ZN(n571) );
  INV_X1 U601 ( .A(n571), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n763) );
  NOR2_X1 U603 ( .A1(n627), .A2(n763), .ZN(n524) );
  XNOR2_X1 U604 ( .A(G128), .B(KEYINPUT29), .ZN(n523) );
  XNOR2_X1 U605 ( .A(n524), .B(n523), .ZN(G30) );
  XNOR2_X1 U606 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n527) );
  XNOR2_X1 U607 ( .A(n526), .B(n527), .ZN(n725) );
  OR2_X1 U608 ( .A1(n725), .A2(n724), .ZN(n728) );
  NOR2_X1 U609 ( .A1(n727), .A2(n728), .ZN(n528) );
  XNOR2_X1 U610 ( .A(n528), .B(KEYINPUT41), .ZN(n741) );
  OR2_X1 U611 ( .A1(n741), .A2(n529), .ZN(n532) );
  INV_X1 U612 ( .A(KEYINPUT115), .ZN(n530) );
  XNOR2_X1 U613 ( .A(n530), .B(KEYINPUT42), .ZN(n531) );
  XNOR2_X1 U614 ( .A(n532), .B(n531), .ZN(n619) );
  XNOR2_X1 U615 ( .A(n619), .B(G137), .ZN(G39) );
  NOR2_X1 U616 ( .A1(n727), .A2(n714), .ZN(n533) );
  XNOR2_X1 U617 ( .A(n533), .B(KEYINPUT108), .ZN(n543) );
  INV_X1 U618 ( .A(G898), .ZN(n536) );
  INV_X1 U619 ( .A(n534), .ZN(n535) );
  NAND2_X1 U620 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U621 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U622 ( .A1(n738), .A2(n539), .ZN(n540) );
  INV_X1 U623 ( .A(n594), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n543), .A2(n569), .ZN(n545) );
  XNOR2_X1 U625 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n544) );
  XNOR2_X1 U626 ( .A(n545), .B(n544), .ZN(n585) );
  NOR2_X1 U627 ( .A1(n362), .A2(n713), .ZN(n547) );
  XNOR2_X1 U628 ( .A(n546), .B(KEYINPUT6), .ZN(n579) );
  NAND2_X1 U629 ( .A1(n547), .A2(n579), .ZN(n548) );
  OR2_X1 U630 ( .A1(n585), .A2(n548), .ZN(n593) );
  XNOR2_X1 U631 ( .A(n593), .B(G101), .ZN(G3) );
  OR2_X1 U632 ( .A1(n550), .A2(n549), .ZN(n760) );
  NOR2_X1 U633 ( .A1(n760), .A2(n551), .ZN(n553) );
  INV_X1 U634 ( .A(n579), .ZN(n552) );
  NAND2_X1 U635 ( .A1(n553), .A2(n552), .ZN(n555) );
  INV_X1 U636 ( .A(KEYINPUT113), .ZN(n554) );
  XNOR2_X1 U637 ( .A(n555), .B(n554), .ZN(n623) );
  INV_X1 U638 ( .A(n623), .ZN(n557) );
  NOR2_X1 U639 ( .A1(n362), .A2(n724), .ZN(n556) );
  NAND2_X1 U640 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U641 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n560), .A2(n526), .ZN(n647) );
  XNOR2_X1 U644 ( .A(n647), .B(G140), .ZN(G42) );
  NOR2_X1 U645 ( .A1(n585), .A2(n362), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n561), .B(KEYINPUT110), .ZN(n563) );
  AND2_X1 U647 ( .A1(n611), .A2(n713), .ZN(n562) );
  XNOR2_X1 U648 ( .A(n587), .B(G110), .ZN(G12) );
  INV_X1 U649 ( .A(KEYINPUT70), .ZN(n565) );
  XNOR2_X2 U650 ( .A(n566), .B(n565), .ZN(n607) );
  XNOR2_X1 U651 ( .A(n595), .B(KEYINPUT111), .ZN(n567) );
  OR2_X2 U652 ( .A1(n567), .A2(n579), .ZN(n568) );
  OR2_X1 U653 ( .A1(n572), .A2(n571), .ZN(n628) );
  XNOR2_X2 U654 ( .A(n573), .B(n382), .ZN(n689) );
  INV_X1 U655 ( .A(KEYINPUT91), .ZN(n574) );
  NAND2_X1 U656 ( .A1(n574), .A2(KEYINPUT44), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n575), .A2(KEYINPUT74), .ZN(n576) );
  INV_X1 U658 ( .A(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n577), .A2(KEYINPUT74), .ZN(n588) );
  INV_X1 U660 ( .A(n588), .ZN(n578) );
  NAND2_X1 U661 ( .A1(n587), .A2(n578), .ZN(n586) );
  XNOR2_X1 U662 ( .A(n579), .B(KEYINPUT83), .ZN(n583) );
  INV_X1 U663 ( .A(n711), .ZN(n581) );
  INV_X1 U664 ( .A(n713), .ZN(n580) );
  OR2_X1 U665 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U666 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n688), .A2(n587), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n604) );
  OR2_X1 U669 ( .A1(KEYINPUT91), .A2(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U670 ( .A1(KEYINPUT74), .A2(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n595), .A2(n546), .ZN(n719) );
  NOR2_X1 U674 ( .A1(n594), .A2(n719), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT31), .ZN(n762) );
  INV_X1 U676 ( .A(n762), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n607), .A2(n608), .ZN(n597) );
  OR2_X1 U678 ( .A1(n597), .A2(n546), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n594), .A2(n598), .ZN(n749) );
  NOR2_X1 U680 ( .A1(n599), .A2(n749), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n763), .B(KEYINPUT106), .ZN(n645) );
  AND2_X1 U682 ( .A1(n645), .A2(n760), .ZN(n729) );
  NOR2_X1 U683 ( .A1(n600), .A2(n729), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U685 ( .A(KEYINPUT88), .B(KEYINPUT45), .Z(n605) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n610) );
  INV_X1 U687 ( .A(n608), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n611), .A2(n724), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT30), .ZN(n613) );
  INV_X1 U691 ( .A(n725), .ZN(n615) );
  INV_X1 U692 ( .A(KEYINPUT75), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT39), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n687), .A2(n619), .ZN(n621) );
  INV_X1 U695 ( .A(KEYINPUT46), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(n643) );
  OR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n625) );
  INV_X1 U698 ( .A(KEYINPUT36), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n625), .B(n624), .ZN(n626) );
  AND2_X1 U700 ( .A1(n626), .A2(n362), .ZN(n765) );
  NOR2_X1 U701 ( .A1(n628), .A2(n526), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n757) );
  NAND2_X1 U703 ( .A1(n632), .A2(KEYINPUT47), .ZN(n634) );
  INV_X1 U704 ( .A(KEYINPUT85), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U706 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n635) );
  NOR2_X1 U707 ( .A1(n729), .A2(n635), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n636), .A2(n627), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  OR2_X1 U711 ( .A1(n646), .A2(n645), .ZN(n686) );
  NAND2_X2 U712 ( .A1(n648), .A2(n424), .ZN(n705) );
  NOR2_X1 U713 ( .A1(n705), .A2(n649), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n767), .A2(n650), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n651), .A2(KEYINPUT2), .ZN(n652) );
  XNOR2_X1 U716 ( .A(n652), .B(KEYINPUT68), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U718 ( .A(n655), .B(KEYINPUT67), .ZN(n657) );
  INV_X1 U719 ( .A(n767), .ZN(n706) );
  NOR2_X2 U720 ( .A1(n657), .A2(n708), .ZN(n692) );
  NAND2_X1 U721 ( .A1(n692), .A2(G475), .ZN(n660) );
  XNOR2_X1 U722 ( .A(n658), .B(KEYINPUT59), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n660), .B(n659), .ZN(n662) );
  INV_X1 U724 ( .A(G952), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n661), .A2(G953), .ZN(n695) );
  NAND2_X1 U726 ( .A1(n662), .A2(n695), .ZN(n664) );
  XOR2_X1 U727 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n663) );
  XNOR2_X1 U728 ( .A(n664), .B(n663), .ZN(G60) );
  NAND2_X1 U729 ( .A1(n692), .A2(G472), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT92), .B(KEYINPUT62), .Z(n665) );
  XNOR2_X1 U731 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n669), .A2(n695), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U735 ( .A1(n692), .A2(G210), .ZN(n675) );
  XNOR2_X1 U736 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT55), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n671), .B(n673), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n695), .ZN(n678) );
  INV_X1 U741 ( .A(KEYINPUT56), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n678), .B(n677), .ZN(G51) );
  NAND2_X1 U743 ( .A1(n692), .A2(G217), .ZN(n681) );
  XOR2_X1 U744 ( .A(n679), .B(KEYINPUT125), .Z(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n682), .A2(n695), .ZN(n684) );
  INV_X1 U747 ( .A(KEYINPUT126), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n684), .B(n683), .ZN(G66) );
  XOR2_X1 U749 ( .A(G134), .B(KEYINPUT119), .Z(n685) );
  XNOR2_X1 U750 ( .A(n686), .B(n685), .ZN(G36) );
  XNOR2_X1 U751 ( .A(n687), .B(G131), .ZN(G33) );
  XNOR2_X1 U752 ( .A(n688), .B(G119), .ZN(G21) );
  BUF_X1 U753 ( .A(n689), .Z(n690) );
  INV_X1 U754 ( .A(n690), .ZN(n691) );
  XOR2_X1 U755 ( .A(n691), .B(G122), .Z(G24) );
  XNOR2_X1 U756 ( .A(n694), .B(n693), .ZN(n696) );
  INV_X1 U757 ( .A(n695), .ZN(n703) );
  NOR2_X1 U758 ( .A1(n696), .A2(n703), .ZN(G63) );
  NAND2_X1 U759 ( .A1(n697), .A2(G469), .ZN(n702) );
  XNOR2_X1 U760 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT58), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(G54) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n707), .A2(KEYINPUT2), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U768 ( .A(n710), .B(KEYINPUT87), .ZN(n746) );
  XOR2_X1 U769 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n722) );
  NOR2_X1 U770 ( .A1(n607), .A2(n362), .ZN(n712) );
  XOR2_X1 U771 ( .A(KEYINPUT50), .B(n712), .Z(n718) );
  NAND2_X1 U772 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U773 ( .A(KEYINPUT49), .B(n715), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n716), .A2(n546), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U777 ( .A(n722), .B(n721), .Z(n723) );
  NOR2_X1 U778 ( .A1(n723), .A2(n741), .ZN(n736) );
  AND2_X1 U779 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U782 ( .A(KEYINPUT121), .B(n730), .Z(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n734) );
  NOR2_X1 U784 ( .A1(n734), .A2(n415), .ZN(n735) );
  NOR2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n737), .B(KEYINPUT52), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n738), .A2(G952), .ZN(n739) );
  NOR2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n744) );
  OR2_X1 U789 ( .A1(n741), .A2(n415), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(n782), .ZN(n743) );
  NOR2_X1 U791 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n746), .A2(n745), .ZN(n748) );
  XOR2_X1 U793 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n747) );
  XNOR2_X1 U794 ( .A(n748), .B(n747), .ZN(G75) );
  INV_X1 U795 ( .A(n749), .ZN(n751) );
  NOR2_X1 U796 ( .A1(n751), .A2(n760), .ZN(n750) );
  XOR2_X1 U797 ( .A(G104), .B(n750), .Z(G6) );
  NOR2_X1 U798 ( .A1(n751), .A2(n763), .ZN(n756) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n753) );
  XNOR2_X1 U800 ( .A(G107), .B(KEYINPUT26), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U802 ( .A(KEYINPUT116), .B(n754), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(G9) );
  XNOR2_X1 U804 ( .A(G143), .B(n757), .ZN(G45) );
  NOR2_X1 U805 ( .A1(n627), .A2(n760), .ZN(n758) );
  XOR2_X1 U806 ( .A(KEYINPUT118), .B(n758), .Z(n759) );
  XNOR2_X1 U807 ( .A(G146), .B(n759), .ZN(G48) );
  NOR2_X1 U808 ( .A1(n760), .A2(n762), .ZN(n761) );
  XOR2_X1 U809 ( .A(G113), .B(n761), .Z(G15) );
  NOR2_X1 U810 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U811 ( .A(G116), .B(n764), .Z(G18) );
  XNOR2_X1 U812 ( .A(n765), .B(G125), .ZN(n766) );
  XNOR2_X1 U813 ( .A(n766), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U814 ( .A1(n767), .A2(n782), .ZN(n771) );
  NAND2_X1 U815 ( .A1(G953), .A2(G224), .ZN(n768) );
  XNOR2_X1 U816 ( .A(KEYINPUT61), .B(n768), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G898), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n771), .A2(n770), .ZN(n776) );
  XOR2_X1 U819 ( .A(n772), .B(G101), .Z(n774) );
  NOR2_X1 U820 ( .A1(n782), .A2(G898), .ZN(n773) );
  NOR2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U822 ( .A(n776), .B(n775), .ZN(G69) );
  XOR2_X1 U823 ( .A(n778), .B(n777), .Z(n779) );
  XNOR2_X1 U824 ( .A(KEYINPUT127), .B(n779), .ZN(n780) );
  XOR2_X1 U825 ( .A(n781), .B(n780), .Z(n784) );
  XNOR2_X1 U826 ( .A(n705), .B(n784), .ZN(n783) );
  NAND2_X1 U827 ( .A1(n783), .A2(n782), .ZN(n788) );
  XNOR2_X1 U828 ( .A(n784), .B(G227), .ZN(n785) );
  NAND2_X1 U829 ( .A1(n785), .A2(G900), .ZN(n786) );
  NAND2_X1 U830 ( .A1(n786), .A2(G953), .ZN(n787) );
  NAND2_X1 U831 ( .A1(n788), .A2(n787), .ZN(G72) );
endmodule

