//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n445, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT72), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(G160));
  AND3_X1   g055(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT73), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT73), .B1(new_n467), .B2(new_n469), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n473), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT74), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n476), .A2(G138), .A3(new_n473), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n473), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G102), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n467), .A2(new_n469), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n473), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n515), .A2(new_n521), .A3(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(G50), .A3(G543), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n519), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n516), .B2(new_n517), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT76), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT77), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT7), .Z(new_n532));
  AOI22_X1  g107(.A1(new_n521), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(new_n514), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(G543), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n532), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(new_n521), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n525), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n541), .A2(new_n548), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT78), .Z(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n536), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n536), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n541), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  INV_X1    g140(.A(G78), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n534), .A2(new_n565), .B1(new_n566), .B2(new_n511), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI221_X1 g144(.A(KEYINPUT79), .B1(new_n566), .B2(new_n511), .C1(new_n534), .C2(new_n565), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(G651), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n562), .A2(new_n564), .A3(new_n571), .ZN(G299));
  XNOR2_X1  g147(.A(G171), .B(KEYINPUT80), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n515), .A2(new_n521), .A3(G87), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n536), .ZN(G288));
  INV_X1    g154(.A(new_n536), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(KEYINPUT83), .A3(G48), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n536), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n581), .A2(new_n584), .B1(new_n563), .B2(G86), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n515), .A2(new_n586), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT81), .B1(new_n534), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(KEYINPUT82), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n591), .B2(G651), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n585), .B1(new_n593), .B2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n580), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n598), .B2(new_n541), .C1(new_n525), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n534), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(KEYINPUT85), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(G651), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n580), .A2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n563), .A2(new_n610), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT84), .B1(new_n541), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT10), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n601), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n601), .B1(G868), .B2(new_n616), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(new_n619), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n551), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT86), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n484), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n487), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  AND2_X1   g213(.A1(new_n473), .A2(G2104), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n476), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT87), .B(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n651), .B(new_n656), .Z(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(G14), .ZN(G401));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(KEYINPUT17), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(new_n662), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n663), .B(KEYINPUT88), .Z(new_n670));
  OAI211_X1 g245(.A(new_n665), .B(new_n669), .C1(new_n667), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT89), .B(G2096), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n676), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n680), .A2(KEYINPUT20), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n676), .A3(new_n679), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n685), .C1(KEYINPUT20), .C2(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1991), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(G229));
  AND2_X1   g268(.A1(KEYINPUT91), .A2(G29), .ZN(new_n694));
  NOR2_X1   g269(.A1(KEYINPUT91), .A2(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT24), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G34), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G160), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G2084), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT31), .B(G11), .ZN(new_n708));
  INV_X1    g283(.A(G171), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G5), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G1961), .ZN(new_n717));
  INV_X1    g292(.A(G1961), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n714), .A2(new_n718), .A3(new_n715), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n551), .A2(new_n711), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n711), .B2(G19), .ZN(new_n721));
  INV_X1    g296(.A(G1341), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n726), .A2(new_n727), .A3(G29), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n723), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  AND4_X1   g304(.A1(new_n708), .A2(new_n717), .A3(new_n719), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G21), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G168), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n697), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n697), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n637), .A2(new_n697), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n711), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n616), .B2(new_n711), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n739), .B1(new_n741), .B2(G1348), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n730), .A2(new_n734), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n492), .A2(new_n696), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n697), .A2(G35), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n744), .A2(KEYINPUT29), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT29), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n746), .A2(new_n747), .B1(KEYINPUT100), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT100), .B(G2090), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G128), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n483), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT96), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G140), .B2(new_n487), .ZN(new_n757));
  OR2_X1    g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G26), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n696), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n697), .A2(KEYINPUT28), .A3(G26), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n711), .A2(G20), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(G29), .A2(G32), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n484), .A2(G129), .B1(G105), .B2(new_n639), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n487), .A2(G141), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(new_n703), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(G29), .A2(G33), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n487), .A2(G139), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n639), .A2(G103), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n785), .B(new_n788), .C1(new_n790), .C2(new_n473), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(new_n703), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n704), .A2(new_n705), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n774), .A2(new_n783), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n741), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n797), .A2(new_n798), .B1(new_n793), .B2(new_n792), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n781), .A2(new_n782), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n768), .A2(new_n796), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n743), .A2(new_n752), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n803));
  NAND2_X1  g378(.A1(G305), .A2(G16), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n711), .A2(G6), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n711), .A2(G23), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G288), .B2(G16), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G1976), .ZN(new_n816));
  AOI211_X1 g391(.A(KEYINPUT33), .B(new_n811), .C1(G288), .C2(G16), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(G1976), .B1(new_n814), .B2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n805), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G305), .B2(G16), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(new_n808), .ZN(new_n824));
  NAND2_X1  g399(.A1(G166), .A2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G1971), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G22), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n711), .B1(new_n524), .B2(new_n528), .ZN(new_n830));
  OAI21_X1  g405(.A(G1971), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n810), .A2(new_n821), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT95), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n808), .A2(new_n823), .B1(new_n829), .B2(new_n831), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n821), .A4(new_n810), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(KEYINPUT34), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n697), .A2(G25), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n484), .A2(G119), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n487), .A2(G131), .ZN(new_n841));
  OR2_X1    g416(.A1(G95), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n839), .B1(new_n845), .B2(new_n697), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G1991), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT92), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n846), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT34), .B1(new_n834), .B2(new_n837), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  MUX2_X1   g427(.A(G24), .B(G290), .S(G16), .Z(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT93), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G1986), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n803), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NOR4_X1   g432(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT36), .A4(new_n855), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n707), .B(new_n802), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(G311));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n852), .A2(new_n803), .A3(new_n856), .ZN(new_n863));
  INV_X1    g438(.A(new_n851), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n864), .A2(new_n856), .A3(new_n838), .A4(new_n849), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT36), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(KEYINPUT102), .A3(new_n707), .A4(new_n802), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n868), .ZN(G150));
  AOI22_X1  g444(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n525), .ZN(new_n871));
  INV_X1    g446(.A(G93), .ZN(new_n872));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  OAI22_X1  g448(.A1(new_n541), .A2(new_n872), .B1(new_n536), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n871), .B2(new_n874), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G860), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n616), .A2(G559), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n551), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n871), .A2(new_n874), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n551), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT104), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(new_n883), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n882), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n879), .B1(new_n890), .B2(G860), .ZN(G145));
  XOR2_X1   g466(.A(new_n492), .B(new_n637), .Z(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n484), .A2(G130), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n487), .A2(G142), .ZN(new_n895));
  OR2_X1    g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n757), .A2(new_n509), .A3(new_n759), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n509), .B1(new_n757), .B2(new_n759), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n760), .A2(G164), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n898), .A3(new_n900), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n791), .B(new_n641), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n909));
  OAI21_X1  g484(.A(G160), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n905), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n702), .A3(new_n907), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n780), .B(new_n844), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n910), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n893), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n914), .ZN(new_n922));
  INV_X1    g497(.A(new_n916), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n892), .A3(new_n917), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n920), .A2(new_n925), .A3(new_n928), .A4(new_n921), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G395));
  XNOR2_X1  g505(.A(G305), .B(G290), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G166), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n931), .A2(G166), .ZN(new_n934));
  OAI21_X1  g509(.A(G288), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  INV_X1    g511(.A(G288), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n889), .A2(new_n626), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n887), .A2(new_n625), .A3(new_n888), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n616), .ZN(new_n944));
  INV_X1    g519(.A(G299), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n616), .A2(KEYINPUT106), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT41), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n943), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT107), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n955), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n940), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n940), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n876), .A2(new_n619), .A3(new_n877), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(G295));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n961), .ZN(G331));
  NOR2_X1   g538(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(G168), .A2(new_n709), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(G301), .B2(G168), .ZN(new_n969));
  INV_X1    g544(.A(new_n888), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT104), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n968), .ZN(new_n973));
  XOR2_X1   g548(.A(G171), .B(KEYINPUT80), .Z(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(G286), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n887), .A2(new_n975), .A3(new_n888), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n954), .A2(new_n952), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n950), .A3(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n938), .B(new_n935), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n976), .ZN(new_n981));
  INV_X1    g556(.A(new_n952), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT41), .B1(new_n948), .B2(new_n949), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n933), .A2(G288), .A3(new_n934), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n937), .B1(new_n936), .B2(new_n932), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n984), .B(new_n978), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n987), .A3(new_n921), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n980), .A2(new_n987), .A3(new_n990), .A4(new_n921), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n964), .B(new_n967), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  AND4_X1   g567(.A1(new_n965), .A2(new_n989), .A3(new_n966), .A4(new_n991), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(KEYINPUT124), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NOR4_X1   g571(.A1(new_n474), .A2(new_n475), .A3(new_n996), .A4(new_n479), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n503), .B2(new_n508), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1001), .A3(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n1005), .B2(new_n737), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  AND4_X1   g583(.A1(KEYINPUT112), .A2(new_n509), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT112), .B1(new_n998), .B2(new_n1007), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n474), .ZN(new_n1012));
  INV_X1    g587(.A(new_n479), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n472), .A2(new_n465), .A3(new_n473), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(G40), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n509), .A2(new_n1008), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1961), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n509), .A2(new_n1008), .A3(new_n999), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n997), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n737), .A2(KEYINPUT53), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT123), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n494), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n495), .A2(new_n500), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G2105), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(KEYINPUT4), .ZN(new_n1028));
  INV_X1    g603(.A(new_n508), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1007), .B(new_n1008), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n998), .A2(KEYINPUT112), .A3(new_n1007), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n997), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n718), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1006), .B1(new_n1024), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n995), .B1(new_n1040), .B2(G301), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  INV_X1    g617(.A(new_n999), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1015), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1004), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n1002), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1046), .B2(G2078), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT124), .A3(new_n974), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1045), .A2(new_n1002), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n477), .A2(new_n478), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n1053), .B(KEYINPUT125), .Z(new_n1054));
  AOI21_X1  g629(.A(new_n996), .B1(new_n1054), .B2(G2105), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1016), .A2(new_n1043), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1047), .B(new_n1036), .C1(new_n1058), .C2(new_n1021), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1059), .A2(new_n974), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1041), .A2(new_n1051), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n937), .A2(G1976), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n998), .A2(G160), .A3(G40), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G288), .A2(new_n816), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1064), .B(new_n1071), .C1(new_n1073), .C2(KEYINPUT52), .ZN(new_n1074));
  INV_X1    g649(.A(G8), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT114), .B(new_n1075), .C1(new_n997), .C2(new_n998), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1068), .B2(G8), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT115), .B(new_n1064), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1072), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1005), .A2(G1971), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT113), .B(G2090), .Z(new_n1088));
  NOR2_X1   g663(.A1(new_n1035), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1086), .B(G8), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n585), .C1(new_n593), .C2(new_n595), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n585), .A2(new_n592), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G1981), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1096), .A3(KEYINPUT49), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1092), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1083), .A2(new_n1090), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n997), .B1(new_n1007), .B2(new_n998), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1030), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1088), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n826), .B2(new_n1046), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1075), .B1(new_n1106), .B2(KEYINPUT116), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1088), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1017), .A2(new_n1030), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1005), .B2(G1971), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1086), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1086), .ZN(new_n1115));
  OAI21_X1  g690(.A(G8), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1106), .A2(KEYINPUT116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1074), .A2(new_n1082), .B1(new_n1092), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1090), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1040), .A2(G301), .B1(new_n1059), .B2(G171), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1017), .A2(new_n1032), .A3(new_n705), .A4(new_n1034), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n733), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G168), .A2(new_n1075), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(G8), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1075), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1128), .B(KEYINPUT121), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT51), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1124), .A2(KEYINPUT54), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT56), .B(G2072), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1044), .B(new_n1141), .C1(new_n1045), .C2(new_n1002), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT57), .B1(new_n945), .B2(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  NAND3_X1  g720(.A1(G299), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n773), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1142), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1068), .A2(G2067), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1035), .B2(new_n798), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n944), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT118), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1152), .A2(KEYINPUT118), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1149), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1996), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1159), .B(new_n1044), .C1(new_n1045), .C2(new_n1002), .ZN(new_n1160));
  OR2_X1    g735(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1161));
  NAND2_X1  g736(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1068), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1160), .A2(KEYINPUT119), .A3(new_n1163), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n551), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1166), .A2(new_n551), .A3(new_n1169), .A4(new_n1167), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n616), .B(new_n1150), .C1(new_n1035), .C2(new_n798), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT60), .B1(new_n1152), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1155), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1149), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1147), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1151), .A2(new_n1181), .A3(new_n616), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1175), .A2(new_n1176), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1158), .B1(new_n1173), .B2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1063), .A2(new_n1123), .A3(new_n1140), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1101), .A2(new_n816), .A3(new_n937), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(new_n1094), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1120), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n1187), .A2(new_n1091), .B1(new_n1188), .B2(new_n1090), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1130), .A2(G286), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1118), .A2(new_n1120), .A3(new_n1090), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(G8), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1194), .B2(new_n1115), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1195), .A2(new_n1120), .A3(new_n1090), .A4(new_n1190), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1189), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1139), .A2(new_n1129), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1198), .A2(new_n1199), .B1(new_n1051), .B2(new_n1041), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1139), .A2(new_n1129), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(KEYINPUT62), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1123), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1185), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1056), .A2(new_n1015), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n760), .B(new_n767), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n780), .B(new_n1159), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n845), .A2(new_n848), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n845), .A2(new_n848), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(G290), .A2(G1986), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1211), .A2(KEYINPUT110), .ZN(new_n1212));
  NAND2_X1  g787(.A1(G290), .A2(G1986), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1212), .B(new_n1213), .Z(new_n1214));
  OAI21_X1  g789(.A(new_n1205), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1204), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1205), .A2(new_n1159), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT46), .Z(new_n1218));
  INV_X1    g793(.A(new_n780), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1206), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1218), .B1(new_n1205), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT47), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1210), .A2(new_n1205), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1205), .A2(new_n1211), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1225), .B(KEYINPUT48), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1228));
  OAI22_X1  g803(.A1(new_n1228), .A2(new_n1208), .B1(G2067), .B2(new_n760), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1229), .A2(new_n1205), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1223), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1223), .A2(KEYINPUT127), .A3(new_n1227), .A4(new_n1230), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1216), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g811(.A1(G227), .A2(G401), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n989), .B2(new_n991), .ZN(new_n1239));
  NOR2_X1   g813(.A1(G229), .A2(new_n463), .ZN(new_n1240));
  NAND3_X1  g814(.A1(new_n926), .A2(new_n1239), .A3(new_n1240), .ZN(G225));
  INV_X1    g815(.A(G225), .ZN(G308));
endmodule


