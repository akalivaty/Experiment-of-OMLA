//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n641, new_n644, new_n646, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(G112), .B2(new_n463), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT67), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n463), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n482), .B(new_n486), .C1(G124), .C2(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n478), .A2(new_n467), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n463), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n479), .B2(new_n480), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n463), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n487), .B2(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n508), .A2(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT68), .B(G51), .Z(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n508), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n511), .A2(new_n510), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n507), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n522), .B2(G64), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n519), .B1(new_n505), .B2(new_n506), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n507), .A2(new_n522), .A3(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n508), .A2(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n522), .A2(G56), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n517), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n511), .A2(new_n510), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT70), .B1(new_n520), .B2(new_n521), .ZN(new_n558));
  OAI21_X1  g133(.A(G65), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n560));
  INV_X1    g135(.A(G78), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n519), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n556), .B1(new_n511), .B2(new_n510), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n520), .A2(KEYINPUT70), .A3(new_n521), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n561), .A2(new_n519), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT71), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n562), .A2(G651), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT69), .ZN(new_n571));
  OAI21_X1  g146(.A(G53), .B1(new_n570), .B2(KEYINPUT69), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n508), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n539), .A2(KEYINPUT69), .A3(new_n570), .A4(G53), .ZN(new_n574));
  INV_X1    g149(.A(new_n514), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n573), .A2(new_n574), .B1(G91), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n569), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G64), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n531), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n579), .B2(new_n536), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(new_n540), .A3(new_n541), .ZN(G301));
  OR2_X1    g156(.A1(new_n530), .A2(new_n534), .ZN(G286));
  NAND2_X1  g157(.A1(new_n539), .A2(G50), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n583), .B1(new_n515), .B2(new_n514), .C1(new_n584), .C2(new_n517), .ZN(G303));
  NOR3_X1   g160(.A1(new_n511), .A2(new_n510), .A3(G74), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT73), .B1(new_n586), .B2(new_n517), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n520), .A2(new_n588), .A3(new_n521), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(new_n590), .A3(G651), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n587), .A2(new_n591), .B1(new_n575), .B2(G87), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n539), .A2(new_n593), .A3(G49), .ZN(new_n594));
  OAI211_X1 g169(.A(G49), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT72), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n539), .A2(KEYINPUT75), .A3(G48), .ZN(new_n599));
  OAI211_X1 g174(.A(G48), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n531), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n599), .A2(new_n602), .B1(new_n605), .B2(G651), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n514), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n507), .A2(new_n522), .A3(KEYINPUT74), .A4(G86), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(G305));
  INV_X1    g186(.A(G60), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n531), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(G72), .A2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g192(.A(KEYINPUT76), .B(G651), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n575), .A2(G85), .B1(G47), .B2(new_n539), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT77), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n617), .A2(new_n622), .A3(new_n618), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n575), .A2(KEYINPUT10), .A3(G92), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n514), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G66), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n564), .B2(new_n565), .ZN(new_n632));
  AND2_X1   g207(.A1(G79), .A2(G543), .ZN(new_n633));
  OAI21_X1  g208(.A(G651), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n539), .A2(G54), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n625), .B1(new_n637), .B2(G868), .ZN(G284));
  OAI21_X1  g213(.A(new_n625), .B1(new_n637), .B2(G868), .ZN(G321));
  NAND2_X1  g214(.A1(G286), .A2(G868), .ZN(new_n640));
  INV_X1    g215(.A(G299), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G868), .ZN(G280));
  XOR2_X1   g217(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n637), .B1(new_n644), .B2(G860), .ZN(G148));
  NOR2_X1   g220(.A1(new_n550), .A2(G868), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n637), .A2(new_n644), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(G868), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g225(.A1(new_n491), .A2(new_n468), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n481), .A2(G135), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n487), .A2(G123), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n463), .A2(G111), .ZN(new_n657));
  OAI21_X1  g232(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(KEYINPUT14), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2451), .B(G2454), .Z(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n669), .B(new_n672), .Z(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  OAI21_X1  g249(.A(G14), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(KEYINPUT81), .A3(new_n674), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(G401));
  XOR2_X1   g255(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT17), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  INV_X1    g263(.A(new_n681), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2096), .B(G2100), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(KEYINPUT20), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n699), .B1(new_n696), .B2(new_n700), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n709), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G6), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G305), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n716), .A2(G23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G288), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G22), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n726), .A2(KEYINPUT85), .A3(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT85), .B1(new_n726), .B2(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(G166), .C2(new_n716), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1971), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n718), .A2(new_n719), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n722), .A2(new_n723), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n725), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT34), .ZN(new_n734));
  MUX2_X1   g309(.A(G24), .B(G290), .S(G16), .Z(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1986), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n481), .A2(G131), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n487), .A2(G119), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n463), .A2(G107), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n741), .S(G29), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT84), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(KEYINPUT86), .B2(KEYINPUT36), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n734), .A2(new_n736), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G34), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(G34), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n751), .B1(new_n753), .B2(KEYINPUT89), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(KEYINPUT89), .B2(new_n753), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G160), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n637), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G4), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n481), .A2(G139), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n764), .B(new_n767), .C1(new_n463), .C2(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G33), .B(new_n769), .S(G29), .Z(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n716), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n716), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n550), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G16), .B2(G19), .ZN(new_n776));
  INV_X1    g351(.A(G1341), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G11), .Z(new_n780));
  INV_X1    g355(.A(G28), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(KEYINPUT30), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT91), .Z(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n781), .B2(KEYINPUT30), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n659), .B2(new_n752), .ZN(new_n786));
  INV_X1    g361(.A(G1961), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n716), .A2(G5), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G301), .B2(G16), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n787), .A2(new_n789), .B1(new_n773), .B2(G1966), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n786), .B(new_n790), .C1(new_n787), .C2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n771), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n762), .B(new_n792), .C1(new_n761), .C2(new_n760), .ZN(new_n793));
  NOR2_X1   g368(.A1(G29), .A2(G35), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G162), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n716), .A2(G20), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT23), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G299), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n752), .A2(G26), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT28), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n481), .A2(G140), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n487), .A2(G128), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n463), .A2(G116), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n806), .B1(new_n811), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT87), .B(G2067), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G27), .A2(G29), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G164), .B2(G29), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n752), .A2(G32), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT26), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n822), .A2(new_n823), .B1(G105), .B2(new_n468), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n481), .A2(G141), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n487), .A2(G129), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n819), .B1(new_n828), .B2(new_n752), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT90), .Z(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT27), .B(G1996), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n814), .B(new_n818), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n797), .A2(new_n798), .ZN(new_n833));
  AOI211_X1 g408(.A(new_n832), .B(new_n833), .C1(new_n831), .C2(new_n830), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n793), .A2(new_n800), .A3(new_n804), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n749), .A2(new_n835), .ZN(G311));
  OR2_X1    g411(.A1(new_n749), .A2(new_n835), .ZN(G150));
  NAND2_X1  g412(.A1(new_n637), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  INV_X1    g415(.A(G80), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n531), .A2(new_n840), .B1(new_n841), .B2(new_n519), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT94), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n844));
  OAI221_X1 g419(.A(new_n844), .B1(new_n841), .B2(new_n519), .C1(new_n531), .C2(new_n840), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(G651), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n575), .A2(G93), .B1(G55), .B2(new_n539), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n549), .B2(new_n546), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n550), .A2(new_n846), .A3(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n839), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n848), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT95), .Z(G145));
  XNOR2_X1  g434(.A(new_n769), .B(new_n828), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n481), .A2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n487), .A2(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n463), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n652), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n769), .B(new_n827), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n811), .B(new_n503), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n741), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n659), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(G162), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n873), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(new_n868), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT96), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n874), .B2(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(G37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(G299), .A2(new_n637), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n569), .A2(new_n636), .A3(new_n576), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT98), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n890));
  AOI211_X1 g465(.A(new_n890), .B(KEYINPUT41), .C1(new_n885), .C2(new_n886), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n851), .B(new_n647), .Z(new_n893));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n636), .B1(new_n569), .B2(new_n576), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n885), .A2(new_n894), .A3(new_n886), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n893), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n893), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  NAND2_X1  g480(.A1(G290), .A2(G288), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n621), .A2(new_n597), .A3(new_n592), .A4(new_n623), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT100), .ZN(new_n909));
  XNOR2_X1  g484(.A(G303), .B(KEYINPUT99), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G305), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n912), .A3(new_n907), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(KEYINPUT101), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n905), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n905), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G868), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n848), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n538), .B2(new_n542), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n580), .A2(KEYINPUT102), .A3(new_n540), .A4(new_n541), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(G168), .ZN(new_n929));
  NOR3_X1   g504(.A1(G171), .A2(G168), .A3(KEYINPUT102), .ZN(new_n930));
  INV_X1    g505(.A(new_n850), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n550), .B1(new_n846), .B2(new_n847), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n929), .A2(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(G286), .A2(G301), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n928), .A3(G168), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n849), .A2(new_n850), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT103), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(KEYINPUT103), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n892), .B2(new_n900), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n936), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n899), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n936), .A2(KEYINPUT103), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n933), .A2(new_n936), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(KEYINPUT103), .ZN(new_n946));
  INV_X1    g521(.A(new_n886), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n888), .B1(new_n947), .B2(new_n896), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n890), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n887), .A2(KEYINPUT98), .A3(new_n888), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  INV_X1    g529(.A(new_n942), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n943), .A2(new_n916), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n892), .A2(new_n900), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n942), .B1(new_n958), .B2(new_n946), .ZN(new_n959));
  INV_X1    g534(.A(new_n916), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT43), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n953), .A3(new_n955), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n941), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n899), .B1(new_n946), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n888), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n916), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND4_X1   g544(.A1(KEYINPUT43), .A2(new_n963), .A3(new_n964), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n957), .B2(new_n961), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n973), .A2(new_n963), .A3(new_n964), .A4(new_n969), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n492), .A2(G2105), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n464), .B2(new_n465), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n980), .A2(KEYINPUT4), .B1(new_n491), .B2(new_n493), .ZN(new_n981));
  OAI211_X1 g556(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n499), .A2(new_n500), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n978), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G125), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n489), .B2(new_n490), .ZN(new_n989));
  INV_X1    g564(.A(new_n474), .ZN(new_n990));
  OAI21_X1  g565(.A(G2105), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(G40), .A3(new_n466), .A4(new_n469), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT124), .Z(new_n998));
  INV_X1    g573(.A(new_n993), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n811), .B(G2067), .Z(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(new_n828), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n996), .B2(new_n995), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT125), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT125), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n827), .B(new_n994), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n741), .A2(new_n744), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n811), .A2(G2067), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n999), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n741), .B(new_n744), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n993), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT126), .Z(new_n1019));
  NOR2_X1   g594(.A1(G290), .A2(G1986), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n993), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1015), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1007), .A2(new_n1009), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n470), .A2(new_n475), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT113), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1029), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n985), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT113), .B1(new_n1035), .B2(new_n1027), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1033), .A2(new_n1036), .A3(G2090), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n992), .B1(new_n985), .B2(new_n986), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1971), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT55), .B(G8), .C1(new_n516), .C2(new_n525), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT106), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT106), .ZN(new_n1044));
  NAND4_X1  g619(.A1(G303), .A2(new_n1044), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(G166), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1027), .B1(new_n985), .B2(new_n1034), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1031), .B1(new_n503), .B2(new_n978), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1049), .C1(new_n1054), .C2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT107), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n987), .A2(new_n1039), .A3(new_n1027), .ZN(new_n1057));
  INV_X1    g632(.A(G1971), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n992), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n798), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(G8), .A4(new_n1049), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n587), .A2(new_n591), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n575), .A2(G87), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n597), .A3(G1976), .A4(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1067), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT109), .B(G1976), .Z(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n592), .B2(new_n597), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT110), .B1(new_n1074), .B2(KEYINPUT52), .ZN(new_n1075));
  INV_X1    g650(.A(new_n591), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n590), .B1(new_n589), .B2(G651), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n597), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1071), .A2(new_n1075), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT75), .B1(new_n539), .B2(G48), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n600), .A2(new_n601), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1086), .A2(new_n1087), .B1(new_n1088), .B2(new_n517), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n609), .A2(new_n610), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(G1981), .ZN(new_n1091));
  INV_X1    g666(.A(G1981), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n514), .A2(new_n608), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n606), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1085), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1047), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1097));
  OAI21_X1  g672(.A(G1981), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n606), .A2(new_n1092), .A3(new_n609), .A4(new_n610), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT49), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT108), .B(new_n1082), .C1(new_n1097), .C2(new_n1070), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1067), .A2(G8), .A3(new_n1070), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(KEYINPUT52), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1084), .B(new_n1101), .C1(new_n1102), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1966), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1057), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1060), .A2(new_n757), .A3(new_n1061), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1047), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(G168), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1051), .A2(new_n1066), .A3(new_n1107), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT114), .B(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1049), .B1(new_n1063), .B2(G8), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1106), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1106), .A2(new_n1119), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1066), .B(new_n1118), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1106), .B(new_n1119), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1066), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G288), .A2(G1976), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1101), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1099), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(KEYINPUT112), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1097), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1128), .B2(KEYINPUT112), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1124), .A2(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1051), .A2(new_n1066), .A3(new_n1107), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1051), .A2(new_n1066), .A3(new_n1107), .A4(KEYINPUT122), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1109), .A2(G168), .A3(new_n1110), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G8), .ZN(new_n1139));
  NAND2_X1  g714(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1138), .A2(G8), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1111), .A2(G286), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT62), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n787), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1038), .A2(KEYINPUT53), .A3(new_n817), .A4(new_n1039), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1057), .B2(G2078), .ZN(new_n1152));
  AOI21_X1  g727(.A(G301), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1139), .A2(new_n1141), .B1(G286), .B2(new_n1111), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1144), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1123), .B(new_n1132), .C1(new_n1137), .C2(new_n1157), .ZN(new_n1158));
  AND4_X1   g733(.A1(G301), .A2(new_n1152), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT54), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1152), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G171), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1150), .A2(G301), .A3(new_n1152), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1160), .A2(new_n1165), .B1(new_n1154), .B2(new_n1144), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1135), .A2(new_n1166), .A3(new_n1136), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n1170));
  XNOR2_X1  g745(.A(G299), .B(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT117), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n641), .A2(new_n1170), .ZN(new_n1174));
  NOR2_X1   g749(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT117), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT115), .B(G1956), .Z(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT56), .B(G2072), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1038), .A2(new_n1039), .A3(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1173), .B(new_n1176), .C1(new_n1181), .C2(KEYINPUT116), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT116), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1067), .A2(G2067), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1187), .B2(new_n761), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n1182), .A2(new_n1185), .B1(new_n636), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1181), .A2(new_n1171), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT58), .B(G1341), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1067), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1192), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1195), .B(new_n1196), .C1(G1996), .C2(new_n1057), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n550), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(KEYINPUT119), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT120), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT59), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1201), .A2(KEYINPUT119), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1197), .A2(new_n1200), .A3(new_n550), .A4(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1188), .A2(KEYINPUT60), .A3(new_n636), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1199), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1181), .A2(new_n1206), .A3(new_n1171), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1171), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1190), .B1(new_n1208), .B2(KEYINPUT61), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1197), .A2(new_n1200), .A3(new_n550), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1188), .A2(KEYINPUT60), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n636), .B1(new_n1188), .B2(KEYINPUT60), .ZN(new_n1212));
  AOI22_X1  g787(.A1(new_n1201), .A2(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1205), .A2(new_n1207), .A3(new_n1209), .A4(new_n1213), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1167), .A2(new_n1168), .B1(new_n1191), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1158), .B1(new_n1169), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1217));
  NAND2_X1  g792(.A1(G290), .A2(G1986), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n999), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1025), .B1(new_n1216), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g795(.A1(G227), .A2(new_n461), .ZN(new_n1222));
  NOR3_X1   g796(.A1(G229), .A2(G401), .A3(new_n1222), .ZN(new_n1223));
  OAI211_X1 g797(.A(new_n883), .B(new_n1223), .C1(new_n974), .C2(new_n975), .ZN(G225));
  INV_X1    g798(.A(G225), .ZN(G308));
endmodule


