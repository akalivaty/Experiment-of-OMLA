

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764;

  AND2_X1 U377 ( .A1(n383), .A2(G472), .ZN(n355) );
  NOR2_X2 U378 ( .A1(n701), .A2(n517), .ZN(n539) );
  AND2_X1 U379 ( .A1(n381), .A2(n379), .ZN(n369) );
  BUF_X1 U380 ( .A(n367), .Z(n368) );
  NAND2_X1 U381 ( .A1(n366), .A2(n633), .ZN(n383) );
  AND2_X1 U382 ( .A1(n528), .A2(n364), .ZN(n372) );
  NOR2_X1 U383 ( .A1(n531), .A2(KEYINPUT45), .ZN(n378) );
  OR2_X1 U384 ( .A1(n716), .A2(n517), .ZN(n390) );
  OR2_X1 U385 ( .A1(n538), .A2(n708), .ZN(n701) );
  INV_X1 U386 ( .A(KEYINPUT64), .ZN(n398) );
  INV_X1 U387 ( .A(n499), .ZN(n356) );
  XNOR2_X1 U388 ( .A(n489), .B(n488), .ZN(n705) );
  BUF_X1 U389 ( .A(n634), .Z(n357) );
  XNOR2_X2 U390 ( .A(n458), .B(n457), .ZN(n751) );
  XNOR2_X2 U391 ( .A(n435), .B(KEYINPUT4), .ZN(n458) );
  XNOR2_X2 U392 ( .A(n498), .B(n669), .ZN(n708) );
  XNOR2_X1 U393 ( .A(G146), .B(G125), .ZN(n424) );
  XNOR2_X1 U394 ( .A(KEYINPUT66), .B(G101), .ZN(n459) );
  XOR2_X1 U395 ( .A(G107), .B(G122), .Z(n436) );
  XOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT105), .Z(n438) );
  XOR2_X1 U397 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n422) );
  XNOR2_X1 U398 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  XNOR2_X1 U399 ( .A(G119), .B(G116), .ZN(n405) );
  XNOR2_X1 U400 ( .A(G137), .B(G140), .ZN(n474) );
  XOR2_X1 U401 ( .A(KEYINPUT12), .B(G140), .Z(n429) );
  XNOR2_X1 U402 ( .A(n751), .B(n460), .ZN(n497) );
  XOR2_X1 U403 ( .A(n549), .B(KEYINPUT86), .Z(n550) );
  AND2_X1 U404 ( .A1(n753), .A2(n621), .ZN(n389) );
  AND2_X1 U405 ( .A1(n753), .A2(n625), .ZN(n388) );
  XNOR2_X1 U406 ( .A(G116), .B(KEYINPUT106), .ZN(n437) );
  XNOR2_X1 U407 ( .A(n423), .B(n391), .ZN(n425) );
  XNOR2_X1 U408 ( .A(KEYINPUT11), .B(KEYINPUT102), .ZN(n421) );
  XNOR2_X1 U409 ( .A(G113), .B(G143), .ZN(n426) );
  INV_X1 U410 ( .A(KEYINPUT95), .ZN(n393) );
  XNOR2_X1 U411 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n395) );
  XNOR2_X1 U412 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U413 ( .A(KEYINPUT77), .B(KEYINPUT91), .Z(n399) );
  INV_X1 U414 ( .A(G902), .ZN(n483) );
  XNOR2_X1 U415 ( .A(G113), .B(KEYINPUT69), .ZN(n404) );
  XNOR2_X1 U416 ( .A(G128), .B(G110), .ZN(n476) );
  XNOR2_X1 U417 ( .A(G110), .B(G107), .ZN(n461) );
  INV_X1 U418 ( .A(G953), .ZN(n699) );
  BUF_X1 U419 ( .A(n716), .Z(n734) );
  OR2_X1 U420 ( .A1(n586), .A2(n571), .ZN(n573) );
  OR2_X1 U421 ( .A1(n670), .A2(G902), .ZN(n498) );
  INV_X1 U422 ( .A(n708), .ZN(n566) );
  XOR2_X1 U423 ( .A(KEYINPUT121), .B(n641), .Z(n642) );
  XNOR2_X1 U424 ( .A(n649), .B(n648), .ZN(n650) );
  OR2_X1 U425 ( .A1(n754), .A2(G952), .ZN(n673) );
  BUF_X1 U426 ( .A(n532), .Z(n763) );
  XNOR2_X1 U427 ( .A(n386), .B(n384), .ZN(G75) );
  XNOR2_X1 U428 ( .A(n385), .B(KEYINPUT120), .ZN(n384) );
  NAND2_X1 U429 ( .A1(n732), .A2(n358), .ZN(n386) );
  INV_X1 U430 ( .A(KEYINPUT53), .ZN(n385) );
  AND2_X1 U431 ( .A1(n731), .A2(n362), .ZN(n358) );
  NOR2_X1 U432 ( .A1(n517), .A2(n542), .ZN(n359) );
  AND2_X1 U433 ( .A1(n499), .A2(n708), .ZN(n360) );
  XOR2_X1 U434 ( .A(n365), .B(KEYINPUT19), .Z(n361) );
  OR2_X1 U435 ( .A1(n734), .A2(n733), .ZN(n362) );
  XOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n363) );
  AND2_X1 U437 ( .A1(n527), .A2(n376), .ZN(n364) );
  NAND2_X1 U438 ( .A1(n561), .A2(n392), .ZN(n365) );
  NAND2_X1 U439 ( .A1(n561), .A2(n392), .ZN(n599) );
  NAND2_X1 U440 ( .A1(n367), .A2(G478), .ZN(n643) );
  BUF_X1 U441 ( .A(n366), .Z(n630) );
  XNOR2_X1 U442 ( .A(n599), .B(KEYINPUT19), .ZN(n581) );
  NAND2_X1 U443 ( .A1(n369), .A2(n377), .ZN(n366) );
  NAND2_X1 U444 ( .A1(n369), .A2(n377), .ZN(n629) );
  NAND2_X1 U445 ( .A1(n628), .A2(n627), .ZN(n371) );
  NAND2_X1 U446 ( .A1(n630), .A2(n753), .ZN(n696) );
  AND2_X2 U447 ( .A1(n371), .A2(n383), .ZN(n367) );
  AND2_X2 U448 ( .A1(n371), .A2(n383), .ZN(n647) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n387) );
  NAND2_X1 U450 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U451 ( .A(n387), .B(n424), .ZN(n397) );
  XNOR2_X2 U452 ( .A(n573), .B(n572), .ZN(n612) );
  XNOR2_X1 U453 ( .A(n370), .B(n577), .ZN(n593) );
  NAND2_X1 U454 ( .A1(n762), .A2(n764), .ZN(n370) );
  AND2_X1 U455 ( .A1(n371), .A2(n355), .ZN(n672) );
  NAND2_X1 U456 ( .A1(n372), .A2(n550), .ZN(n381) );
  NAND2_X1 U457 ( .A1(n375), .A2(n373), .ZN(n377) );
  NAND2_X1 U458 ( .A1(n550), .A2(n374), .ZN(n373) );
  INV_X1 U459 ( .A(n378), .ZN(n374) );
  OR2_X1 U460 ( .A1(n550), .A2(KEYINPUT45), .ZN(n375) );
  NAND2_X1 U461 ( .A1(n528), .A2(n527), .ZN(n382) );
  INV_X1 U462 ( .A(KEYINPUT45), .ZN(n376) );
  NAND2_X1 U463 ( .A1(n382), .A2(n380), .ZN(n379) );
  AND2_X1 U464 ( .A1(n531), .A2(KEYINPUT45), .ZN(n380) );
  NAND2_X1 U465 ( .A1(n368), .A2(G217), .ZN(n662) );
  NAND2_X1 U466 ( .A1(n368), .A2(G469), .ZN(n667) );
  NAND2_X1 U467 ( .A1(n383), .A2(n698), .ZN(n700) );
  NAND2_X1 U468 ( .A1(n366), .A2(n388), .ZN(n626) );
  NAND2_X1 U469 ( .A1(n629), .A2(n389), .ZN(n622) );
  INV_X1 U470 ( .A(n616), .ZN(n617) );
  AND2_X1 U471 ( .A1(G214), .A2(n490), .ZN(n391) );
  NAND2_X1 U472 ( .A1(n414), .A2(G214), .ZN(n392) );
  INV_X1 U473 ( .A(KEYINPUT110), .ZN(n469) );
  XNOR2_X1 U474 ( .A(n425), .B(n472), .ZN(n432) );
  BUF_X1 U475 ( .A(n540), .Z(n565) );
  XNOR2_X1 U476 ( .A(n434), .B(n433), .ZN(n534) );
  INV_X1 U477 ( .A(KEYINPUT122), .ZN(n645) );
  XNOR2_X1 U478 ( .A(n576), .B(n575), .ZN(n762) );
  XNOR2_X2 U479 ( .A(KEYINPUT94), .B(KEYINPUT17), .ZN(n394) );
  XNOR2_X1 U480 ( .A(n459), .B(n395), .ZN(n396) );
  XNOR2_X1 U481 ( .A(n397), .B(n396), .ZN(n403) );
  XNOR2_X2 U482 ( .A(n398), .B(G953), .ZN(n462) );
  NAND2_X1 U483 ( .A1(n462), .A2(G224), .ZN(n400) );
  XNOR2_X2 U484 ( .A(G143), .B(G128), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n401), .B(n458), .ZN(n402) );
  XNOR2_X1 U486 ( .A(n403), .B(n402), .ZN(n410) );
  XNOR2_X1 U487 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U488 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U489 ( .A(n407), .B(n406), .ZN(n495) );
  XNOR2_X1 U490 ( .A(G104), .B(G122), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n428), .B(KEYINPUT16), .ZN(n408) );
  XNOR2_X1 U492 ( .A(n408), .B(n461), .ZN(n409) );
  XNOR2_X1 U493 ( .A(n495), .B(n409), .ZN(n743) );
  XNOR2_X1 U494 ( .A(n410), .B(n743), .ZN(n634) );
  NAND2_X1 U495 ( .A1(n634), .A2(n623), .ZN(n413) );
  INV_X1 U496 ( .A(G237), .ZN(n411) );
  NAND2_X1 U497 ( .A1(n483), .A2(n411), .ZN(n414) );
  AND2_X1 U498 ( .A1(n414), .A2(G210), .ZN(n412) );
  XNOR2_X2 U499 ( .A(n413), .B(n412), .ZN(n561) );
  NOR2_X1 U500 ( .A1(G898), .A2(n699), .ZN(n744) );
  NAND2_X1 U501 ( .A1(n744), .A2(G902), .ZN(n415) );
  NAND2_X1 U502 ( .A1(n699), .A2(G952), .ZN(n552) );
  NAND2_X1 U503 ( .A1(n415), .A2(n552), .ZN(n418) );
  NAND2_X1 U504 ( .A1(G237), .A2(G234), .ZN(n417) );
  INV_X1 U505 ( .A(KEYINPUT14), .ZN(n416) );
  XNOR2_X1 U506 ( .A(n417), .B(n416), .ZN(n729) );
  INV_X1 U507 ( .A(n729), .ZN(n554) );
  AND2_X1 U508 ( .A1(n418), .A2(n554), .ZN(n419) );
  NAND2_X1 U509 ( .A1(n581), .A2(n419), .ZN(n420) );
  XNOR2_X1 U510 ( .A(n420), .B(KEYINPUT0), .ZN(n516) );
  XNOR2_X1 U511 ( .A(n422), .B(n421), .ZN(n423) );
  NOR2_X1 U512 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U513 ( .A(KEYINPUT10), .B(n424), .ZN(n472) );
  XNOR2_X1 U514 ( .A(G131), .B(n426), .ZN(n427) );
  XNOR2_X1 U515 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U516 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U517 ( .A(n432), .B(n431), .ZN(n649) );
  NAND2_X1 U518 ( .A1(n649), .A2(n483), .ZN(n434) );
  XNOR2_X1 U519 ( .A(KEYINPUT13), .B(G475), .ZN(n433) );
  XNOR2_X1 U520 ( .A(n435), .B(n436), .ZN(n440) );
  XNOR2_X1 U521 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U522 ( .A(n440), .B(n439), .Z(n443) );
  NAND2_X1 U523 ( .A1(n462), .A2(G234), .ZN(n441) );
  XOR2_X1 U524 ( .A(KEYINPUT8), .B(n441), .Z(n471) );
  NAND2_X1 U525 ( .A1(G217), .A2(n471), .ZN(n442) );
  XNOR2_X1 U526 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U527 ( .A(G134), .B(KEYINPUT9), .Z(n444) );
  XNOR2_X1 U528 ( .A(n445), .B(n444), .ZN(n641) );
  NAND2_X1 U529 ( .A1(n641), .A2(n483), .ZN(n447) );
  XNOR2_X1 U530 ( .A(KEYINPUT107), .B(G478), .ZN(n446) );
  XNOR2_X1 U531 ( .A(n447), .B(n446), .ZN(n535) );
  NAND2_X1 U532 ( .A1(n534), .A2(n535), .ZN(n719) );
  XOR2_X1 U533 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n449) );
  NAND2_X1 U534 ( .A1(G234), .A2(n623), .ZN(n448) );
  XNOR2_X1 U535 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U536 ( .A(KEYINPUT98), .B(n450), .ZN(n484) );
  NAND2_X1 U537 ( .A1(G221), .A2(n484), .ZN(n452) );
  XOR2_X1 U538 ( .A(KEYINPUT21), .B(KEYINPUT100), .Z(n451) );
  XNOR2_X1 U539 ( .A(n452), .B(n451), .ZN(n706) );
  INV_X1 U540 ( .A(n706), .ZN(n453) );
  OR2_X1 U541 ( .A1(n719), .A2(n453), .ZN(n454) );
  NOR2_X2 U542 ( .A1(n516), .A2(n454), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n455), .B(n363), .ZN(n503) );
  INV_X1 U544 ( .A(G131), .ZN(n456) );
  XNOR2_X1 U545 ( .A(n456), .B(G134), .ZN(n457) );
  XNOR2_X1 U546 ( .A(n459), .B(G146), .ZN(n460) );
  XNOR2_X1 U547 ( .A(KEYINPUT96), .B(n474), .ZN(n748) );
  XNOR2_X1 U548 ( .A(n461), .B(G104), .ZN(n464) );
  BUF_X2 U549 ( .A(n462), .Z(n754) );
  NAND2_X1 U550 ( .A1(n754), .A2(G227), .ZN(n463) );
  XNOR2_X1 U551 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U552 ( .A(n748), .B(n465), .ZN(n466) );
  XNOR2_X1 U553 ( .A(n497), .B(n466), .ZN(n665) );
  OR2_X2 U554 ( .A1(n665), .A2(G902), .ZN(n467) );
  XNOR2_X2 U555 ( .A(n467), .B(G469), .ZN(n540) );
  INV_X1 U556 ( .A(KEYINPUT1), .ZN(n468) );
  XNOR2_X2 U557 ( .A(n540), .B(n468), .ZN(n703) );
  NAND2_X1 U558 ( .A1(n503), .A2(n703), .ZN(n470) );
  XNOR2_X1 U559 ( .A(n470), .B(n469), .ZN(n500) );
  NAND2_X1 U560 ( .A1(G221), .A2(n471), .ZN(n473) );
  INV_X1 U561 ( .A(n472), .ZN(n749) );
  XNOR2_X1 U562 ( .A(n473), .B(n749), .ZN(n482) );
  INV_X1 U563 ( .A(n474), .ZN(n475) );
  XNOR2_X1 U564 ( .A(n476), .B(n475), .ZN(n480) );
  XOR2_X1 U565 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n478) );
  XNOR2_X1 U566 ( .A(G119), .B(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U567 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U568 ( .A(n480), .B(n479), .Z(n481) );
  XNOR2_X1 U569 ( .A(n482), .B(n481), .ZN(n661) );
  NAND2_X1 U570 ( .A1(n661), .A2(n483), .ZN(n489) );
  NAND2_X1 U571 ( .A1(G217), .A2(n484), .ZN(n487) );
  INV_X1 U572 ( .A(KEYINPUT76), .ZN(n485) );
  XNOR2_X1 U573 ( .A(n485), .B(KEYINPUT25), .ZN(n486) );
  XNOR2_X1 U574 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U575 ( .A(n705), .ZN(n499) );
  NAND2_X1 U576 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n491), .B(G137), .ZN(n493) );
  XNOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT5), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U580 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U581 ( .A(n497), .B(n496), .ZN(n670) );
  INV_X1 U582 ( .A(G472), .ZN(n669) );
  NAND2_X1 U583 ( .A1(n500), .A2(n360), .ZN(n502) );
  INV_X1 U584 ( .A(KEYINPUT111), .ZN(n501) );
  XNOR2_X1 U585 ( .A(n502), .B(n501), .ZN(n677) );
  BUF_X1 U586 ( .A(n503), .Z(n504) );
  XNOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT6), .ZN(n505) );
  XNOR2_X1 U588 ( .A(n708), .B(n505), .ZN(n596) );
  XNOR2_X1 U589 ( .A(n596), .B(KEYINPUT79), .ZN(n507) );
  OR2_X1 U590 ( .A1(n703), .A2(n356), .ZN(n506) );
  NOR2_X1 U591 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U592 ( .A1(n504), .A2(n508), .ZN(n509) );
  XNOR2_X1 U593 ( .A(n509), .B(KEYINPUT32), .ZN(n660) );
  NAND2_X1 U594 ( .A1(n677), .A2(n660), .ZN(n511) );
  INV_X1 U595 ( .A(KEYINPUT88), .ZN(n510) );
  XNOR2_X2 U596 ( .A(n511), .B(n510), .ZN(n530) );
  NOR2_X1 U597 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n512) );
  XNOR2_X1 U598 ( .A(n530), .B(n512), .ZN(n526) );
  NAND2_X1 U599 ( .A1(n705), .A2(n706), .ZN(n702) );
  NOR2_X1 U600 ( .A1(n703), .A2(n702), .ZN(n513) );
  XNOR2_X1 U601 ( .A(n513), .B(KEYINPUT75), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n538), .A2(n596), .ZN(n515) );
  XNOR2_X1 U603 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n514) );
  XNOR2_X1 U604 ( .A(n515), .B(n514), .ZN(n716) );
  BUF_X1 U605 ( .A(n516), .Z(n517) );
  XOR2_X1 U606 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n518) );
  XNOR2_X1 U607 ( .A(n390), .B(n518), .ZN(n520) );
  OR2_X1 U608 ( .A1(n535), .A2(n534), .ZN(n587) );
  INV_X1 U609 ( .A(n587), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n523) );
  INV_X1 U611 ( .A(KEYINPUT83), .ZN(n521) );
  XNOR2_X1 U612 ( .A(n521), .B(KEYINPUT35), .ZN(n522) );
  XNOR2_X1 U613 ( .A(n523), .B(n522), .ZN(n532) );
  INV_X1 U614 ( .A(KEYINPUT44), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n763), .A2(n524), .ZN(n525) );
  INV_X1 U616 ( .A(KEYINPUT65), .ZN(n527) );
  NAND2_X1 U617 ( .A1(KEYINPUT44), .A2(KEYINPUT65), .ZN(n529) );
  OR2_X1 U618 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U619 ( .A1(n532), .A2(KEYINPUT44), .ZN(n548) );
  INV_X1 U620 ( .A(n535), .ZN(n533) );
  AND2_X1 U621 ( .A1(n533), .A2(n534), .ZN(n692) );
  INV_X1 U622 ( .A(n534), .ZN(n536) );
  AND2_X1 U623 ( .A1(n536), .A2(n535), .ZN(n690) );
  NOR2_X1 U624 ( .A1(n692), .A2(n690), .ZN(n537) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT108), .ZN(n720) );
  XNOR2_X1 U626 ( .A(KEYINPUT80), .B(n720), .ZN(n579) );
  XOR2_X1 U627 ( .A(n539), .B(KEYINPUT31), .Z(n693) );
  NOR2_X1 U628 ( .A1(n566), .A2(n702), .ZN(n541) );
  NAND2_X1 U629 ( .A1(n541), .A2(n565), .ZN(n542) );
  NOR2_X1 U630 ( .A1(n693), .A2(n359), .ZN(n543) );
  NOR2_X1 U631 ( .A1(n579), .A2(n543), .ZN(n546) );
  AND2_X1 U632 ( .A1(n596), .A2(n356), .ZN(n544) );
  AND2_X1 U633 ( .A1(n544), .A2(n703), .ZN(n545) );
  AND2_X1 U634 ( .A1(n504), .A2(n545), .ZN(n680) );
  NOR2_X1 U635 ( .A1(n546), .A2(n680), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U637 ( .A1(G900), .A2(n754), .ZN(n551) );
  NAND2_X1 U638 ( .A1(G902), .A2(n551), .ZN(n553) );
  NAND2_X1 U639 ( .A1(n553), .A2(n552), .ZN(n555) );
  AND2_X1 U640 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U641 ( .A1(n706), .A2(n556), .ZN(n564) );
  INV_X1 U642 ( .A(n564), .ZN(n557) );
  OR2_X1 U643 ( .A1(n705), .A2(n557), .ZN(n594) );
  OR2_X1 U644 ( .A1(n594), .A2(n708), .ZN(n559) );
  INV_X1 U645 ( .A(KEYINPUT28), .ZN(n558) );
  XNOR2_X1 U646 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U647 ( .A1(n560), .A2(n565), .ZN(n582) );
  BUF_X1 U648 ( .A(n561), .Z(n616) );
  XNOR2_X1 U649 ( .A(n616), .B(KEYINPUT38), .ZN(n571) );
  INV_X1 U650 ( .A(n571), .ZN(n717) );
  NAND2_X1 U651 ( .A1(n717), .A2(n392), .ZN(n721) );
  NOR2_X1 U652 ( .A1(n719), .A2(n721), .ZN(n562) );
  XNOR2_X1 U653 ( .A(KEYINPUT41), .B(n562), .ZN(n733) );
  OR2_X1 U654 ( .A1(n582), .A2(n733), .ZN(n563) );
  XNOR2_X1 U655 ( .A(n563), .B(KEYINPUT42), .ZN(n764) );
  NAND2_X1 U656 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n566), .A2(n392), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n567), .B(KEYINPUT30), .ZN(n568) );
  NOR2_X1 U659 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n570), .A2(n356), .ZN(n586) );
  XOR2_X1 U661 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n572) );
  NAND2_X1 U662 ( .A1(n612), .A2(n690), .ZN(n576) );
  XOR2_X1 U663 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n574) );
  XNOR2_X1 U664 ( .A(KEYINPUT40), .B(n574), .ZN(n575) );
  XNOR2_X1 U665 ( .A(KEYINPUT85), .B(KEYINPUT46), .ZN(n577) );
  XOR2_X1 U666 ( .A(KEYINPUT67), .B(KEYINPUT47), .Z(n578) );
  NOR2_X1 U667 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U668 ( .A(n580), .B(KEYINPUT74), .ZN(n583) );
  NOR2_X1 U669 ( .A1(n582), .A2(n361), .ZN(n687) );
  AND2_X1 U670 ( .A1(n583), .A2(n687), .ZN(n591) );
  INV_X1 U671 ( .A(n720), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n584), .A2(n687), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n585), .A2(KEYINPUT47), .ZN(n589) );
  NOR2_X1 U674 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n616), .A2(n588), .ZN(n655) );
  NAND2_X1 U676 ( .A1(n589), .A2(n655), .ZN(n590) );
  NOR2_X1 U677 ( .A1(n591), .A2(n590), .ZN(n592) );
  AND2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n607) );
  INV_X1 U679 ( .A(n594), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n690), .A2(n595), .ZN(n597) );
  OR2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT112), .ZN(n614) );
  XNOR2_X1 U683 ( .A(n614), .B(KEYINPUT115), .ZN(n601) );
  INV_X1 U684 ( .A(n365), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n603) );
  XNOR2_X1 U686 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n603), .B(n602), .ZN(n605) );
  INV_X1 U688 ( .A(n703), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U690 ( .A(n606), .B(KEYINPUT116), .ZN(n659) );
  NAND2_X1 U691 ( .A1(n607), .A2(n659), .ZN(n611) );
  XNOR2_X1 U692 ( .A(KEYINPUT84), .B(KEYINPUT48), .ZN(n609) );
  INV_X1 U693 ( .A(KEYINPUT68), .ZN(n608) );
  XNOR2_X1 U694 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U695 ( .A(n611), .B(n610), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n612), .A2(n692), .ZN(n695) );
  NAND2_X1 U697 ( .A1(n703), .A2(n392), .ZN(n613) );
  OR2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n615), .B(KEYINPUT43), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n656) );
  AND2_X1 U701 ( .A1(n695), .A2(n656), .ZN(n619) );
  AND2_X2 U702 ( .A1(n620), .A2(n619), .ZN(n753) );
  INV_X1 U703 ( .A(KEYINPUT81), .ZN(n621) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n697) );
  NAND2_X1 U705 ( .A1(n622), .A2(n697), .ZN(n624) );
  INV_X1 U706 ( .A(n623), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n624), .A2(n625), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n626), .A2(KEYINPUT81), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n753), .A2(KEYINPUT2), .ZN(n632) );
  INV_X1 U710 ( .A(KEYINPUT82), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n647), .A2(G210), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n635) );
  XNOR2_X1 U714 ( .A(n357), .B(n635), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n638), .A2(n673), .ZN(n640) );
  INV_X1 U717 ( .A(KEYINPUT56), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n640), .B(n639), .ZN(G51) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n644), .A2(n673), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(G63) );
  NAND2_X1 U722 ( .A1(n647), .A2(G475), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT92), .B(KEYINPUT59), .Z(n648) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n673), .ZN(n654) );
  INV_X1 U726 ( .A(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G60) );
  XNOR2_X1 U728 ( .A(n655), .B(G143), .ZN(G45) );
  XNOR2_X1 U729 ( .A(n656), .B(G140), .ZN(G42) );
  XOR2_X1 U730 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n657) );
  XOR2_X1 U731 ( .A(n657), .B(G125), .Z(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(G27) );
  XNOR2_X1 U733 ( .A(n660), .B(G119), .ZN(G21) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  AND2_X1 U735 ( .A1(n663), .A2(n673), .ZN(G66) );
  XNOR2_X1 U736 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(n668) );
  AND2_X1 U739 ( .A1(n668), .A2(n673), .ZN(G54) );
  XNOR2_X1 U740 ( .A(n670), .B(KEYINPUT62), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U743 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G57) );
  BUF_X1 U745 ( .A(n677), .Z(n678) );
  XOR2_X1 U746 ( .A(G110), .B(KEYINPUT117), .Z(n679) );
  XNOR2_X1 U747 ( .A(n678), .B(n679), .ZN(G12) );
  XOR2_X1 U748 ( .A(G101), .B(n680), .Z(G3) );
  NAND2_X1 U749 ( .A1(n359), .A2(n690), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(G104), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U752 ( .A1(n359), .A2(n692), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U754 ( .A(G107), .B(n684), .ZN(G9) );
  XOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  NAND2_X1 U756 ( .A1(n687), .A2(n692), .ZN(n685) );
  XNOR2_X1 U757 ( .A(n686), .B(n685), .ZN(G30) );
  NAND2_X1 U758 ( .A1(n687), .A2(n690), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT118), .ZN(n689) );
  XNOR2_X1 U760 ( .A(G146), .B(n689), .ZN(G48) );
  NAND2_X1 U761 ( .A1(n693), .A2(n690), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n691), .B(G113), .ZN(G15) );
  NAND2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(G116), .ZN(G18) );
  XNOR2_X1 U765 ( .A(G134), .B(n695), .ZN(G36) );
  NAND2_X1 U766 ( .A1(n696), .A2(n697), .ZN(n698) );
  AND2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n732) );
  INV_X1 U768 ( .A(n701), .ZN(n713) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U770 ( .A(KEYINPUT50), .B(n704), .Z(n711) );
  NOR2_X1 U771 ( .A1(n706), .A2(n356), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT49), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U776 ( .A(KEYINPUT51), .B(n714), .Z(n715) );
  NOR2_X1 U777 ( .A1(n733), .A2(n715), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n717), .A2(n392), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U781 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n734), .A2(n724), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n727), .B(KEYINPUT52), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U786 ( .A1(G952), .A2(n730), .ZN(n731) );
  INV_X1 U787 ( .A(n630), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n735), .A2(G953), .ZN(n741) );
  XOR2_X1 U789 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n737) );
  NAND2_X1 U790 ( .A1(G224), .A2(G953), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U792 ( .A1(G898), .A2(n738), .ZN(n739) );
  XOR2_X1 U793 ( .A(KEYINPUT124), .B(n739), .Z(n740) );
  NOR2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT125), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n743), .B(G101), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(G69) );
  XOR2_X1 U799 ( .A(KEYINPUT126), .B(n748), .Z(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n756) );
  XOR2_X1 U802 ( .A(n753), .B(n756), .Z(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n761) );
  XNOR2_X1 U804 ( .A(G227), .B(n756), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(G900), .ZN(n758) );
  XOR2_X1 U806 ( .A(KEYINPUT127), .B(n758), .Z(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(n759), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(G72) );
  XNOR2_X1 U809 ( .A(G131), .B(n762), .ZN(G33) );
  XOR2_X1 U810 ( .A(n763), .B(G122), .Z(G24) );
  XNOR2_X1 U811 ( .A(G137), .B(n764), .ZN(G39) );
endmodule

