//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(G50gat), .B(G78gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n208), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G141gat), .B(G148gat), .Z(new_n214));
  AOI22_X1  g013(.A1(new_n214), .A2(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n210), .B(KEYINPUT73), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218));
  INV_X1    g017(.A(G211gat), .ZN(new_n219));
  INV_X1    g018(.A(G218gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G211gat), .B(G218gat), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT29), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n226), .B(new_n227), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n234));
  AOI21_X1  g033(.A(new_n217), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n226), .A2(new_n227), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n209), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n214), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n209), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n210), .B(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n239), .B(new_n234), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n207), .B1(new_n235), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n245), .A2(KEYINPUT81), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(KEYINPUT81), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n237), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n207), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n206), .B1(new_n248), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT82), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n205), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n257), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n244), .B1(new_n228), .B2(KEYINPUT80), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(new_n237), .B2(KEYINPUT80), .ZN(new_n263));
  INV_X1    g062(.A(new_n234), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n251), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n256), .B1(new_n265), .B2(new_n246), .ZN(new_n266));
  OAI21_X1  g065(.A(G22gat), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n206), .A3(new_n257), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n267), .A2(new_n259), .A3(new_n268), .A4(new_n205), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  INV_X1    g072(.A(G64gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT23), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n283), .A2(new_n288), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n281), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n288), .A4(new_n290), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n302), .B(new_n303), .C1(new_n284), .C2(new_n285), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT28), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT68), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n306), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT28), .B1(new_n307), .B2(new_n305), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n280), .B(new_n304), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n301), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n278), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n280), .ZN(new_n320));
  INV_X1    g119(.A(new_n306), .ZN(new_n321));
  INV_X1    g120(.A(new_n311), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n322), .A2(new_n323), .A3(new_n308), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT68), .B1(new_n310), .B2(new_n311), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n314), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n320), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n328), .A2(new_n304), .B1(new_n296), .B2(new_n300), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT71), .B(new_n317), .C1(new_n329), .C2(KEYINPUT29), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n315), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n296), .A2(new_n300), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n317), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n232), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n296), .A2(new_n334), .A3(new_n300), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n334), .B1(new_n296), .B2(new_n300), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n315), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n329), .A2(new_n318), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n237), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n277), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT30), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n232), .B1(new_n343), .B2(new_n344), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n341), .A2(new_n318), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n319), .A3(new_n330), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n232), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT72), .B(new_n350), .C1(new_n354), .C2(new_n277), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  INV_X1    g159(.A(G134gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G127gat), .A2(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT69), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G113gat), .ZN(new_n370));
  INV_X1    g169(.A(G113gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G120gat), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT1), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(G120gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n369), .A2(G113gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n362), .A2(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n251), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n217), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n359), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n380), .B(new_n243), .C1(new_n217), .C2(new_n249), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n216), .B(new_n209), .C1(KEYINPUT2), .C2(new_n208), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n389), .A3(new_n390), .A4(new_n239), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n217), .B2(new_n382), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n385), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(KEYINPUT77), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT4), .B1(new_n380), .B2(new_n251), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n217), .A2(new_n398), .A3(new_n390), .A4(new_n382), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n358), .A2(new_n386), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n388), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n402), .A3(new_n408), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n403), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n354), .A2(new_n277), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n356), .A2(new_n357), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n349), .A2(new_n355), .A3(new_n416), .ZN(new_n418));
  INV_X1    g217(.A(new_n415), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT78), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n272), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n272), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT38), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n277), .C1(new_n354), .C2(KEYINPUT37), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n352), .A2(new_n237), .A3(new_n319), .A4(new_n330), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n343), .A2(new_n232), .A3(new_n344), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT37), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT83), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n277), .B1(new_n354), .B2(KEYINPUT37), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n338), .A2(new_n346), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT37), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT38), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n277), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n423), .A4(new_n427), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n415), .A2(new_n347), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n429), .A2(new_n434), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n385), .B1(new_n400), .B2(new_n388), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n384), .A2(new_n386), .ZN(new_n443));
  OR3_X1    g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n409), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT40), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n448), .A3(new_n410), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n422), .B1(new_n440), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n421), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n336), .A2(new_n380), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n341), .A2(new_n382), .ZN(new_n453));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n454), .B(KEYINPUT64), .Z(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G43gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n455), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n336), .A2(new_n380), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n341), .A2(new_n382), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n453), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n456), .A2(KEYINPUT32), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n467), .B2(new_n470), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n470), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n468), .B2(new_n463), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT32), .B(new_n456), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n462), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT36), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  INV_X1    g281(.A(new_n480), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n478), .B2(new_n472), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n451), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n272), .A2(new_n475), .A3(new_n480), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n418), .A2(new_n419), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n272), .A2(new_n475), .A3(new_n480), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n417), .B2(new_n420), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n492), .B2(new_n488), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  OR3_X1    g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n498), .A2(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT15), .A3(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  AOI21_X1  g307(.A(G1gat), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n509), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT86), .B(G8gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT87), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n509), .B(new_n511), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n515), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(new_n513), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n506), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n502), .A2(KEYINPUT17), .A3(new_n504), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT17), .B1(new_n502), .B2(new_n504), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n524), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT88), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT18), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n529), .B(KEYINPUT89), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT13), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT87), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n536), .A2(new_n537), .A3(new_n505), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n538), .B2(new_n524), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n505), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n526), .A2(new_n527), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n522), .A3(new_n520), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n529), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(KEYINPUT88), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n533), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G169gat), .B(G197gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n533), .A2(new_n539), .A3(new_n545), .A4(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n285), .ZN(new_n559));
  INV_X1    g358(.A(G204gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n276), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n565), .B2(new_n276), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G57gat), .B(G64gat), .Z(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  INV_X1    g374(.A(G71gat), .ZN(new_n576));
  INV_X1    g375(.A(G78gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n574), .A2(new_n580), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT90), .B1(new_n582), .B2(new_n583), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n573), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT10), .B(new_n572), .C1(new_n586), .C2(new_n587), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n563), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT10), .B1(new_n588), .B2(new_n589), .ZN(new_n597));
  INV_X1    g396(.A(new_n593), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n595), .B(new_n562), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n588), .A2(new_n563), .A3(new_n589), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n561), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n594), .A2(new_n603), .A3(new_n561), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n557), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n495), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n219), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n536), .A2(new_n537), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n586), .A2(new_n587), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G183gat), .ZN(new_n616));
  INV_X1    g415(.A(G183gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n611), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n616), .B2(new_n618), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n610), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n624), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n624), .B2(new_n628), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n541), .A2(new_n573), .ZN(new_n635));
  AND2_X1   g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n505), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n636), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n305), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G218gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n638), .A2(new_n641), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n642), .B2(new_n646), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n608), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n419), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  INV_X1    g453(.A(new_n418), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n508), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n662), .B(new_n663), .C1(new_n658), .C2(new_n656), .ZN(G1325gat));
  NOR2_X1   g463(.A1(new_n483), .A2(new_n484), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n652), .B2(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT36), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT36), .B1(new_n475), .B2(new_n480), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT94), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT94), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n485), .A2(new_n670), .A3(new_n481), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n651), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n666), .B1(G15gat), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n651), .A2(new_n272), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  OAI21_X1  g476(.A(new_n649), .B1(new_n486), .B2(new_n494), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n634), .A2(new_n607), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G29gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n419), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(new_n649), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n669), .B(new_n671), .C1(new_n421), .C2(new_n450), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT95), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n688), .A2(new_n689), .A3(new_n493), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n688), .B2(new_n493), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT96), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n687), .C1(new_n690), .C2(new_n691), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n697), .A2(new_n419), .A3(new_n680), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n685), .B1(new_n683), .B2(new_n698), .ZN(G1328gat));
  NOR3_X1   g498(.A1(new_n681), .A2(G36gat), .A3(new_n655), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT46), .ZN(new_n701));
  INV_X1    g500(.A(G36gat), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n697), .A2(new_n418), .A3(new_n680), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(G1329gat));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  INV_X1    g504(.A(new_n672), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n697), .A2(new_n706), .A3(new_n680), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT97), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n697), .A2(new_n709), .A3(new_n706), .A4(new_n680), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(G43gat), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(G43gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n682), .A2(new_n712), .A3(new_n665), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n705), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n707), .A2(G43gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n705), .A3(new_n713), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT98), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n719));
  INV_X1    g518(.A(new_n713), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n712), .B1(new_n707), .B2(KEYINPUT97), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n710), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n719), .B(new_n716), .C1(new_n722), .C2(new_n705), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n718), .A2(new_n723), .ZN(G1330gat));
  NAND3_X1  g523(.A1(new_n697), .A2(new_n422), .A3(new_n680), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n681), .A2(G50gat), .A3(new_n272), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT48), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n728), .B(new_n730), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n690), .A2(new_n691), .ZN(new_n732));
  INV_X1    g531(.A(new_n606), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n634), .A2(new_n649), .A3(new_n556), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n419), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g538(.A(new_n655), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT100), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT101), .Z(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1333gat));
  NAND3_X1  g544(.A1(new_n737), .A2(new_n576), .A3(new_n665), .ZN(new_n746));
  OAI21_X1  g545(.A(G71gat), .B1(new_n736), .B2(new_n672), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g548(.A1(new_n736), .A2(new_n272), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n577), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n688), .A2(new_n493), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n634), .A2(new_n557), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n686), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT51), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n757), .A2(new_n606), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n419), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n754), .A2(new_n733), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n697), .A2(G85gat), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n419), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n697), .A2(new_n418), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n655), .A2(G92gat), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n760), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT102), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(KEYINPUT51), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n753), .A2(new_n756), .A3(new_n771), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n770), .B(KEYINPUT51), .C1(new_n752), .C2(new_n755), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n606), .B(new_n767), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n766), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT103), .B1(new_n775), .B2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g575(.A(new_n774), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n765), .B2(G92gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n769), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT104), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n784), .B(new_n769), .C1(new_n776), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n697), .A2(new_n706), .A3(new_n762), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(G99gat), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n760), .A2(new_n792), .A3(new_n665), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n697), .A2(new_n422), .A3(new_n762), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n733), .A2(G106gat), .A3(new_n272), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n772), .B2(new_n773), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n795), .B2(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n757), .A2(new_n759), .A3(new_n797), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n801), .A2(KEYINPUT106), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT106), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1339gat));
  NAND3_X1  g604(.A1(new_n592), .A2(new_n563), .A3(new_n593), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n594), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n592), .A2(KEYINPUT107), .A3(new_n563), .A4(new_n593), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT54), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n596), .B2(new_n600), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n812), .A3(new_n561), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT55), .A4(new_n561), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n556), .A2(new_n815), .A3(new_n605), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n538), .A2(new_n524), .A3(new_n535), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n529), .B1(new_n540), .B2(new_n542), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n551), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT108), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(new_n551), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(new_n555), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n606), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n649), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n815), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n649), .A2(new_n555), .A3(new_n823), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n816), .A2(new_n605), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n634), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n634), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n686), .A3(new_n733), .A4(new_n557), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT109), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n487), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n419), .A3(new_n655), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n557), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(new_n371), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n840), .B2(new_n733), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n606), .A2(new_n369), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT110), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n840), .B2(new_n845), .ZN(G1341gat));
  OR2_X1    g645(.A1(new_n840), .A2(new_n634), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n847), .A2(new_n848), .A3(new_n360), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(new_n360), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n360), .B2(new_n847), .ZN(G1342gat));
  OAI21_X1  g651(.A(G134gat), .B1(new_n840), .B2(new_n686), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT113), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n686), .A2(new_n418), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT112), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n839), .A2(new_n361), .A3(new_n419), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n859));
  NOR2_X1   g658(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n854), .B(new_n861), .C1(new_n859), .C2(new_n858), .ZN(G1343gat));
  XNOR2_X1  g661(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n813), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n556), .A2(new_n864), .A3(new_n605), .A4(new_n816), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n649), .B1(new_n865), .B2(new_n825), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n634), .B1(new_n866), .B2(new_n830), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n272), .B1(new_n867), .B2(new_n833), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n838), .A2(new_n422), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n706), .A2(new_n415), .A3(new_n418), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n556), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n556), .A4(new_n874), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(G141gat), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n871), .A2(new_n415), .A3(new_n706), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n655), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n557), .A2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n875), .A2(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n886), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT118), .B1(new_n889), .B2(KEYINPUT58), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n891), .B(new_n880), .C1(new_n888), .C2(new_n886), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(G1344gat));
  INV_X1    g692(.A(G148gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n894), .A3(new_n606), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n874), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n733), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n894), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n422), .A4(new_n837), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n634), .A2(new_n649), .A3(new_n606), .A4(new_n556), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n865), .A2(new_n825), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n686), .ZN(new_n906));
  INV_X1    g705(.A(new_n830), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(new_n634), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT120), .B(new_n903), .C1(new_n909), .C2(new_n272), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n900), .A2(new_n902), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n733), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n874), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n896), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n895), .B1(new_n899), .B2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n882), .B2(new_n832), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n897), .A2(new_n634), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(G155gat), .B2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n897), .B2(new_n686), .ZN(new_n920));
  INV_X1    g719(.A(G162gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n881), .A2(new_n921), .A3(new_n857), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n655), .A2(new_n419), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n839), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n557), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(new_n284), .ZN(G1348gat));
  NOR2_X1   g726(.A1(new_n925), .A2(new_n733), .ZN(new_n928));
  XOR2_X1   g727(.A(KEYINPUT121), .B(G176gat), .Z(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1349gat));
  OR4_X1    g729(.A1(new_n634), .A2(new_n925), .A3(new_n325), .A4(new_n324), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n617), .B1(new_n925), .B2(new_n634), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1350gat));
  NOR2_X1   g736(.A1(new_n925), .A2(new_n686), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n305), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT61), .B(G190gat), .Z(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n938), .B2(new_n941), .ZN(G1351gat));
  NAND2_X1  g741(.A1(new_n672), .A2(new_n924), .ZN(new_n943));
  NOR4_X1   g742(.A1(new_n871), .A2(G197gat), .A3(new_n557), .A4(new_n943), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT123), .Z(new_n945));
  NOR2_X1   g744(.A1(new_n912), .A2(new_n943), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n557), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1352gat));
  NOR2_X1   g748(.A1(new_n871), .A2(new_n943), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n560), .A3(new_n606), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  INV_X1    g751(.A(new_n943), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n560), .B1(new_n913), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n911), .A2(new_n832), .A3(new_n953), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n956), .A2(new_n959), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n956), .A2(G211gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n965), .B(KEYINPUT63), .C1(new_n956), .C2(G211gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n219), .A3(new_n832), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n964), .A2(new_n966), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n971), .B(new_n968), .C1(new_n972), .C2(new_n961), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n973), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n947), .B2(new_n686), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n950), .A2(new_n220), .A3(new_n649), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


