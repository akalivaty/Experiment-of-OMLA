//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G57gat), .B(G64gat), .Z(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n202), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n214), .B(new_n215), .Z(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G211gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G8gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(G8gat), .B1(new_n225), .B2(KEYINPUT85), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n212), .A2(new_n213), .ZN(new_n234));
  OAI21_X1  g033(.A(G183gat), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n228), .A2(new_n236), .A3(new_n237), .A4(new_n232), .ZN(new_n238));
  INV_X1    g037(.A(G231gat), .ZN(new_n239));
  INV_X1    g038(.A(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n235), .B2(new_n238), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n220), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n243), .A2(new_n244), .A3(new_n220), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n217), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n216), .A3(new_n245), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT0), .B(G57gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G85gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  XNOR2_X1  g056(.A(G155gat), .B(G162gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260));
  XNOR2_X1  g059(.A(G141gat), .B(G148gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n259), .B(new_n260), .C1(KEYINPUT2), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G141gat), .ZN(new_n264));
  INV_X1    g063(.A(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G148gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT2), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT73), .B1(new_n267), .B2(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n266), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT2), .B1(new_n271), .B2(KEYINPUT74), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n258), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G127gat), .B(G134gat), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(G113gat), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(G113gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G113gat), .B2(new_n279), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n276), .B(new_n277), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G120gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n275), .B1(KEYINPUT1), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n257), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n283), .A2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(new_n273), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(new_n262), .B2(new_n268), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT4), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n269), .A2(new_n294), .A3(new_n273), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n290), .A2(new_n294), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n290), .A2(new_n294), .B1(new_n285), .B2(new_n283), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT75), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n292), .B(new_n293), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n290), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n286), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT5), .B1(new_n307), .B2(new_n293), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n303), .A2(KEYINPUT76), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n303), .B2(KEYINPUT76), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n256), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n312));
  INV_X1    g111(.A(new_n308), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n303), .A2(KEYINPUT76), .A3(new_n308), .ZN(new_n315));
  INV_X1    g114(.A(new_n256), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n309), .A2(new_n310), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT6), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  NOR2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  AND2_X1   g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT24), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n326), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n340), .A2(G169gat), .A3(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .A3(new_n342), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n324), .B1(new_n338), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT64), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n332), .A2(KEYINPUT64), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n337), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT25), .B1(new_n341), .B2(KEYINPUT65), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT65), .B1(new_n325), .B2(KEYINPUT23), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n326), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n352), .A2(new_n342), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  AND2_X1   g156(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT28), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n357), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n325), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n342), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n361), .A2(new_n364), .A3(new_n368), .A4(new_n327), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n323), .B1(new_n348), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n327), .A2(KEYINPUT67), .A3(new_n328), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT67), .B1(new_n327), .B2(new_n328), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n337), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n326), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n344), .A4(new_n346), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT25), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n369), .A3(new_n356), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n372), .B(KEYINPUT71), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n371), .A2(new_n372), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G211gat), .A2(G218gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n388), .A2(new_n389), .B1(new_n390), .B2(new_n383), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT70), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(new_n389), .ZN(new_n395));
  OAI22_X1  g194(.A1(KEYINPUT22), .A2(new_n384), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT70), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT72), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT72), .ZN(new_n401));
  INV_X1    g200(.A(new_n372), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n371), .A2(new_n380), .B1(new_n379), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n403), .B2(new_n399), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n379), .B2(new_n323), .ZN(new_n405));
  INV_X1    g204(.A(new_n370), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n380), .B1(new_n406), .B2(new_n378), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n405), .A2(new_n407), .A3(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n400), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G8gat), .B(G36gat), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G64gat), .ZN(new_n411));
  INV_X1    g210(.A(G92gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n400), .B(new_n413), .C1(new_n404), .C2(new_n408), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT30), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(new_n418), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n322), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n290), .B2(new_n294), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n399), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n393), .A2(new_n397), .A3(new_n323), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n290), .B1(new_n424), .B2(new_n294), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n295), .A2(new_n323), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT78), .A3(new_n398), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n422), .B2(new_n399), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n394), .A2(new_n396), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n391), .A2(new_n386), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n323), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n274), .B1(KEYINPUT3), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT77), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT77), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n274), .B(new_n437), .C1(KEYINPUT3), .C2(new_n434), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n429), .A2(new_n431), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n427), .B1(new_n439), .B2(new_n426), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G22gat), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n443));
  XOR2_X1   g242(.A(G78gat), .B(G106gat), .Z(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n443), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n440), .B2(KEYINPUT79), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n440), .B2(KEYINPUT79), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n421), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n379), .A2(new_n288), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n406), .A2(new_n286), .A3(new_n378), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n456), .A2(new_n457), .A3(G227gat), .A4(G233gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n458), .B(KEYINPUT32), .C1(new_n460), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n456), .A2(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n471), .B(KEYINPUT34), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n465), .A3(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT69), .B1(new_n465), .B2(new_n467), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(new_n475), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n454), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n409), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n371), .A2(new_n372), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n379), .A2(new_n381), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n399), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n401), .C1(new_n399), .C2(new_n403), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(KEYINPUT37), .A3(new_n400), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n413), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT38), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n319), .A3(new_n321), .A4(new_n415), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT81), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n382), .B2(new_n399), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n403), .A2(new_n399), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT81), .B(new_n398), .C1(new_n405), .C2(new_n407), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT38), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n486), .A2(new_n500), .A3(new_n501), .A4(new_n413), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n414), .B1(new_n409), .B2(new_n485), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n501), .A4(new_n500), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n484), .B1(new_n494), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n307), .A2(new_n293), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n287), .A2(new_n291), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT75), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT39), .B(new_n509), .C1(new_n513), .C2(new_n293), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n513), .A2(new_n293), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n256), .B(new_n514), .C1(new_n515), .C2(KEYINPUT39), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n416), .A2(KEYINPUT30), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n413), .B1(new_n490), .B2(new_n400), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n419), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n417), .A2(KEYINPUT80), .A3(new_n419), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n320), .A2(new_n316), .B1(new_n516), .B2(new_n517), .ZN(new_n526));
  AND4_X1   g325(.A1(new_n518), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n455), .B(new_n483), .C1(new_n508), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n525), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n449), .A2(new_n477), .A3(new_n453), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n322), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n454), .A2(new_n482), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n319), .A2(new_n321), .B1(new_n419), .B2(new_n417), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G190gat), .B(G218gat), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT91), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT88), .B(KEYINPUT92), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n545), .A2(new_n546), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(KEYINPUT15), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(KEYINPUT15), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(KEYINPUT15), .A3(new_n548), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(KEYINPUT15), .B2(new_n548), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT7), .ZN(new_n559));
  NAND2_X1  g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  AOI22_X1  g360(.A1(KEYINPUT8), .A2(new_n560), .B1(new_n561), .B2(new_n412), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n557), .A2(KEYINPUT89), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT89), .B1(new_n557), .B2(new_n566), .ZN(new_n568));
  AND2_X1   g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n563), .B(new_n564), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n551), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n567), .A2(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n537), .A2(KEYINPUT91), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n575), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n541), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n578), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n540), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n551), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n233), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n228), .A2(new_n552), .A3(new_n556), .A4(new_n232), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT86), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT18), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n228), .A2(new_n232), .A3(new_n551), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n593), .B(KEYINPUT13), .Z(new_n600));
  NAND3_X1  g399(.A1(new_n233), .A2(KEYINPUT87), .A3(new_n590), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT18), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(KEYINPUT86), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT11), .B(G169gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G197gat), .ZN(new_n607));
  XOR2_X1   g406(.A(G113gat), .B(G141gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT83), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n596), .A2(new_n611), .A3(new_n602), .A4(new_n604), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G230gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n240), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT93), .B1(new_n559), .B2(new_n562), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n571), .B1(new_n212), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n212), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n566), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n566), .A2(new_n621), .A3(KEYINPUT10), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n618), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n618), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT94), .ZN(new_n634));
  INV_X1    g433(.A(G176gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n628), .A2(new_n630), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n616), .A2(new_n640), .ZN(new_n641));
  AND4_X1   g440(.A1(new_n252), .A2(new_n536), .A3(new_n589), .A4(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n322), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT95), .B(G1gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1324gat));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(KEYINPUT97), .A2(KEYINPUT42), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n529), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n651), .B(KEYINPUT96), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(G8gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n642), .B2(new_n477), .ZN(new_n658));
  INV_X1    g457(.A(new_n483), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n642), .A2(G15gat), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n642), .A2(new_n454), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT98), .B(KEYINPUT43), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n447), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n662), .B(new_n664), .ZN(G1327gat));
  AOI21_X1  g464(.A(new_n589), .B1(new_n528), .B2(new_n535), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n641), .A2(new_n251), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(G29gat), .A3(new_n322), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n483), .B1(new_n508), .B2(new_n527), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n421), .A2(KEYINPUT100), .A3(new_n454), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n534), .B2(new_n484), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n535), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n588), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n679), .A2(new_n680), .B1(new_n681), .B2(new_n666), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n668), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n643), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n672), .B1(new_n686), .B2(new_n543), .ZN(G1328gat));
  NOR3_X1   g486(.A1(new_n669), .A2(G36gat), .A3(new_n529), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n684), .A2(new_n650), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n544), .ZN(G1329gat));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n683), .B2(new_n483), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n682), .A2(KEYINPUT103), .A3(new_n659), .A4(new_n668), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(G43gat), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n669), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n478), .A2(G43gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n684), .B2(new_n659), .ZN(new_n704));
  INV_X1    g503(.A(new_n700), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(G1330gat));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n524), .A2(new_n518), .A3(new_n525), .A4(new_n526), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n709), .B(new_n484), .C1(new_n494), .C2(new_n507), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n710), .A2(new_n483), .A3(new_n676), .A4(new_n674), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n589), .B(new_n680), .C1(new_n711), .C2(new_n535), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n681), .B1(new_n536), .B2(new_n588), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n454), .B(new_n668), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(G50gat), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n669), .A2(G50gat), .A3(new_n484), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n708), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n682), .A2(new_n719), .A3(new_n454), .A4(new_n668), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n720), .A3(G50gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n716), .A2(new_n708), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n717), .B1(new_n724), .B2(new_n725), .ZN(G1331gat));
  NOR3_X1   g525(.A1(new_n251), .A2(new_n588), .A3(new_n615), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n678), .A2(new_n640), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n678), .A2(KEYINPUT106), .A3(new_n640), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n643), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n650), .A2(KEYINPUT107), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n529), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  OAI21_X1  g544(.A(new_n205), .B1(new_n732), .B2(new_n478), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n730), .A2(G71gat), .A3(new_n659), .A4(new_n731), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT50), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n753), .B(new_n746), .C1(new_n749), .C2(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1334gat));
  NOR2_X1   g554(.A1(new_n732), .A2(new_n484), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n206), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n252), .A2(new_n615), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n640), .B(new_n758), .C1(new_n712), .C2(new_n713), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n759), .A2(KEYINPUT109), .A3(new_n322), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT109), .B1(new_n759), .B2(new_n322), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(G85gat), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n589), .B1(new_n711), .B2(new_n535), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n758), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n679), .A2(KEYINPUT110), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n766), .A4(new_n758), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n767), .A2(new_n768), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n640), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n643), .A2(new_n561), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n762), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n739), .A2(new_n412), .A3(new_n640), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT112), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n773), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  OAI21_X1  g582(.A(G92gat), .B1(new_n759), .B2(new_n740), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n759), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n412), .B1(new_n786), .B2(new_n650), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n780), .B1(new_n769), .B2(new_n772), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n759), .B2(new_n483), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n478), .A2(G99gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n776), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g592(.A(new_n640), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n484), .A2(G106gat), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT114), .Z(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n773), .A2(new_n775), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND2_X1  g598(.A1(KEYINPUT113), .A2(G106gat), .ZN(new_n800));
  OR2_X1    g599(.A1(KEYINPUT113), .A2(G106gat), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n800), .B(new_n801), .C1(new_n759), .C2(new_n484), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n796), .B1(new_n769), .B2(new_n772), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n616), .A2(G113gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NOR4_X1   g608(.A1(new_n251), .A2(new_n588), .A3(new_n640), .A4(new_n615), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n636), .B1(new_n627), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n625), .A2(new_n618), .A3(new_n626), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n812), .B(KEYINPUT55), .C1(new_n627), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n639), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n639), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n593), .B1(new_n591), .B2(new_n592), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n609), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n614), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n812), .B1(new_n627), .B2(new_n814), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n588), .A2(new_n820), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n824), .A2(new_n794), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n613), .A2(new_n614), .B1(new_n827), .B2(new_n826), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n820), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n832), .B2(new_n588), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n810), .B1(new_n833), .B2(new_n251), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n454), .A2(new_n482), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n809), .B1(new_n837), .B2(new_n643), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n322), .A4(new_n836), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n740), .B(new_n808), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n834), .A2(new_n454), .A3(new_n478), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n739), .A2(new_n322), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n615), .A3(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(KEYINPUT116), .A3(G113gat), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT116), .B1(new_n843), .B2(G113gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(G1340gat));
  NOR2_X1   g647(.A1(new_n838), .A2(new_n839), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n739), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n279), .A3(new_n640), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n841), .A2(new_n842), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852), .B2(new_n794), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n850), .B2(new_n252), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n852), .A2(new_n251), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(G127gat), .B2(new_n856), .ZN(G1342gat));
  INV_X1    g656(.A(new_n849), .ZN(new_n858));
  INV_X1    g657(.A(G134gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n650), .A2(new_n589), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n852), .B2(new_n589), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n833), .A2(new_n251), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(new_n454), .C1(new_n867), .C2(new_n810), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n736), .A2(new_n643), .A3(new_n483), .A4(new_n738), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n816), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n830), .B1(new_n831), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n829), .B1(new_n873), .B2(new_n588), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n810), .B1(new_n874), .B2(new_n251), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n484), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n868), .A2(new_n871), .A3(KEYINPUT120), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n265), .B1(new_n881), .B2(new_n615), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n834), .A2(new_n484), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n643), .A3(new_n483), .ZN(new_n884));
  NOR4_X1   g683(.A1(new_n884), .A2(G141gat), .A3(new_n616), .A4(new_n739), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(G141gat), .B1(new_n877), .B2(new_n616), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n884), .A2(new_n739), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n263), .A3(new_n640), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n263), .C1(new_n881), .C2(new_n640), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n874), .A2(new_n251), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n866), .B(new_n454), .C1(new_n895), .C2(new_n810), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n834), .B2(new_n484), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n871), .A3(new_n640), .A4(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n263), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n894), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n893), .B2(new_n902), .ZN(G1345gat));
  AOI21_X1  g702(.A(G155gat), .B1(new_n891), .B2(new_n252), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n252), .A2(G155gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT122), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n881), .B2(new_n906), .ZN(G1346gat));
  INV_X1    g706(.A(new_n884), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT74), .B(G162gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n860), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n589), .B1(new_n879), .B2(new_n880), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n834), .A2(new_n643), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n739), .A2(KEYINPUT123), .A3(new_n835), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n740), .B2(new_n836), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n917), .A2(G169gat), .A3(new_n616), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n643), .A2(new_n529), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n841), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n616), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(G1348gat));
  INV_X1    g721(.A(new_n917), .ZN(new_n923));
  AOI21_X1  g722(.A(G176gat), .B1(new_n923), .B2(new_n640), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n920), .A2(new_n635), .A3(new_n794), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n252), .A3(new_n362), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  OAI21_X1  g728(.A(G183gat), .B1(new_n920), .B2(new_n251), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n931), .B(new_n932), .Z(G1350gat));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n357), .A3(new_n588), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n920), .B2(new_n589), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  AND2_X1   g737(.A1(new_n896), .A2(new_n897), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n919), .A2(new_n483), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n616), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n834), .A2(new_n643), .A3(new_n659), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n740), .A2(new_n484), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n616), .B2(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n943), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n949), .B2(new_n794), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n949), .A2(KEYINPUT62), .A3(new_n794), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n939), .A2(new_n640), .A3(new_n940), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n948), .ZN(G1353gat));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n896), .A2(new_n897), .A3(new_n252), .A4(new_n940), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n954), .B(KEYINPUT63), .C1(new_n957), .C2(new_n219), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n955), .B(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n959), .A2(G211gat), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n943), .A2(new_n219), .A3(new_n252), .A4(new_n945), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT125), .Z(new_n964));
  NAND3_X1  g763(.A1(new_n958), .A2(new_n962), .A3(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n941), .B2(new_n589), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n589), .A2(G218gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n943), .A2(new_n945), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1355gat));
endmodule


