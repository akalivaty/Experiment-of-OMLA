//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n195), .B2(G146), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n195), .A2(new_n197), .A3(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(G237), .A2(G953), .ZN(new_n202));
  AOI21_X1  g016(.A(G143), .B1(new_n202), .B2(G214), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT18), .A2(G131), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n205), .ZN(new_n208));
  OAI211_X1 g022(.A(KEYINPUT18), .B(G131), .C1(new_n208), .C2(new_n203), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n201), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT19), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT19), .B1(new_n192), .B2(new_n194), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT16), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n208), .B2(new_n203), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n204), .A2(new_n220), .A3(new_n205), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n190), .B1(new_n210), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n201), .A2(new_n207), .A3(new_n209), .ZN(new_n224));
  INV_X1    g038(.A(new_n217), .ZN(new_n225));
  AOI21_X1  g039(.A(G146), .B1(new_n215), .B2(new_n216), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT17), .B(G131), .C1(new_n208), .C2(new_n203), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT87), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n227), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n224), .B(new_n189), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(G475), .A2(G902), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT20), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n224), .B1(new_n232), .B2(new_n233), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(new_n189), .ZN(new_n243));
  OAI21_X1  g057(.A(G475), .B1(new_n243), .B2(G902), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G952), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G953), .ZN(new_n247));
  INV_X1    g061(.A(G234), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT92), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT21), .B(G898), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT93), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n254), .B(new_n255), .C1(G234), .C2(G237), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT88), .B1(new_n259), .B2(G116), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G122), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT14), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n264), .A2(KEYINPUT14), .ZN(new_n268));
  OAI21_X1  g082(.A(G107), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G128), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G143), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT64), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n274), .A3(new_n270), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT64), .B(G134), .ZN(new_n284));
  INV_X1    g098(.A(new_n282), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n275), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n264), .A2(new_n288), .A3(new_n266), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n269), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n264), .A2(new_n266), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G107), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n289), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n273), .B2(G143), .ZN(new_n295));
  INV_X1    g109(.A(new_n272), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT89), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT89), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n271), .A2(G128), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n298), .B(new_n272), .C1(new_n299), .C2(new_n294), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(KEYINPUT13), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n293), .B(new_n286), .C1(new_n302), .C2(new_n277), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  INV_X1    g119(.A(G217), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n305), .A2(new_n306), .A3(G953), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n290), .A2(new_n303), .A3(new_n307), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G478), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n290), .A2(new_n303), .A3(new_n307), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n307), .B1(new_n290), .B2(new_n303), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n254), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n245), .A2(new_n258), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n188), .A2(G107), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n288), .A2(KEYINPUT3), .A3(G104), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT3), .B1(new_n288), .B2(G104), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G101), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n188), .B2(G107), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n288), .A2(KEYINPUT3), .A3(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT79), .A3(new_n333), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n339), .A2(new_n340), .B1(new_n188), .B2(G107), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n333), .B1(new_n345), .B2(new_n337), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n332), .A2(G101), .ZN(new_n347));
  INV_X1    g161(.A(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G116), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n262), .A2(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT2), .B(G113), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n351), .ZN(new_n354));
  INV_X1    g168(.A(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n346), .A2(new_n347), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n288), .B2(G104), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n288), .A2(G104), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n188), .A2(KEYINPUT80), .A3(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G101), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n337), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT81), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n366), .A3(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n369), .A2(G113), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(new_n354), .B2(new_n355), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n344), .A2(new_n357), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G122), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n328), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n373), .B2(KEYINPUT86), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n346), .A2(new_n347), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n356), .A2(new_n353), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT79), .B1(new_n342), .B2(new_n333), .ZN(new_n380));
  NOR4_X1   g194(.A1(new_n345), .A2(new_n335), .A3(KEYINPUT4), .A4(new_n337), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n372), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n375), .B1(new_n377), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n374), .B1(new_n384), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n373), .A2(KEYINPUT86), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n328), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G143), .B(G146), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT0), .A3(G128), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G128), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G125), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT1), .B1(new_n271), .B2(G146), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n271), .A2(G146), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n211), .A2(G143), .ZN(new_n398));
  OAI211_X1 g212(.A(G128), .B(new_n396), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n211), .A2(G143), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n271), .A2(G146), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n400), .B(new_n401), .C1(KEYINPUT1), .C2(new_n273), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n395), .B1(new_n404), .B2(G125), .ZN(new_n405));
  INV_X1    g219(.A(G224), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n387), .A2(new_n390), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n384), .A2(new_n376), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n405), .B1(new_n411), .B2(new_n407), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n407), .A2(new_n411), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n395), .B(new_n413), .C1(new_n404), .C2(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n368), .B(new_n372), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n374), .B(KEYINPUT8), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n409), .A2(new_n420), .A3(new_n422), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n327), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n325), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n255), .A2(G227), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT78), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n399), .A2(KEYINPUT66), .A3(new_n402), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT66), .B1(new_n399), .B2(new_n402), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT10), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n362), .A2(new_n366), .A3(G101), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n366), .B1(new_n362), .B2(G101), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n364), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT82), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n403), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n399), .A2(KEYINPUT66), .A3(new_n402), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n368), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  INV_X1    g262(.A(G137), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(G134), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(G137), .B1(new_n278), .B2(new_n280), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n448), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n281), .A2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n279), .A2(G134), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n277), .A2(KEYINPUT64), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n448), .B(new_n449), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(G131), .B1(new_n284), .B2(G137), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n368), .A2(new_n404), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n394), .B1(new_n346), .B2(new_n347), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n464), .A2(new_n440), .B1(new_n344), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n447), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n447), .B2(new_n466), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT84), .B(new_n432), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n447), .A2(new_n463), .A3(new_n466), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n365), .A2(new_n403), .A3(new_n367), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n403), .B1(new_n365), .B2(new_n367), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT12), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n432), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n435), .A2(new_n438), .A3(KEYINPUT82), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n445), .B1(new_n444), .B2(new_n368), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n466), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n470), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT84), .B1(new_n485), .B2(new_n432), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n428), .B(new_n254), .C1(new_n480), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n470), .A2(new_n478), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n470), .A2(new_n477), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n489), .A2(new_n484), .B1(new_n490), .B2(new_n432), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n488), .B(G469), .C1(new_n491), .C2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n432), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n478), .A3(new_n470), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G469), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n428), .A2(new_n254), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G221), .ZN(new_n500));
  INV_X1    g314(.A(new_n305), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n254), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(KEYINPUT85), .A3(new_n503), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n427), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n500), .A2(new_n248), .A3(G953), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n348), .B2(G128), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n273), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(new_n515), .C1(G119), .C2(new_n273), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n516), .A2(G110), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT74), .ZN(new_n518));
  XNOR2_X1  g332(.A(G119), .B(G128), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT24), .B(G110), .Z(new_n520));
  OAI22_X1  g334(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n518), .B2(new_n517), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n217), .B1(new_n199), .B2(new_n200), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n227), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n516), .A2(G110), .B1(new_n519), .B2(new_n520), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n512), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n511), .C1(new_n522), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n254), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g346(.A1(G217), .A2(G902), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n306), .B2(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT73), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n529), .A2(new_n536), .A3(new_n254), .A4(new_n530), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n529), .A2(new_n530), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n535), .A2(G902), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT76), .Z(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n545));
  NOR2_X1   g359(.A1(G472), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n379), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n449), .A2(G134), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n451), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n220), .B1(new_n281), .B2(new_n449), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n452), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT65), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT65), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n554), .B(new_n550), .C1(new_n452), .C2(new_n551), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(new_n404), .ZN(new_n556));
  INV_X1    g370(.A(new_n394), .ZN(new_n557));
  INV_X1    g371(.A(new_n453), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n220), .B1(new_n459), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n452), .A2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n548), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n552), .B1(new_n443), .B2(new_n442), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n394), .B1(new_n454), .B2(new_n461), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(new_n379), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT28), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n461), .B(new_n550), .C1(new_n433), .C2(new_n434), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n548), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT68), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(KEYINPUT68), .A3(new_n569), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n202), .A2(G210), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n568), .A2(new_n578), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT30), .B1(new_n556), .B2(new_n561), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n442), .A2(new_n443), .ZN(new_n583));
  INV_X1    g397(.A(new_n549), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n284), .B2(G137), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n459), .A2(new_n460), .B1(G131), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n462), .A2(new_n557), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n548), .B1(new_n587), .B2(KEYINPUT30), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n580), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT31), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n574), .A2(new_n579), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n579), .B1(new_n587), .B2(new_n548), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n561), .A2(KEYINPUT30), .A3(new_n567), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n379), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n594), .B2(new_n581), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT67), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT67), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n592), .B(new_n597), .C1(new_n594), .C2(new_n581), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(KEYINPUT31), .A3(new_n598), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n545), .B(new_n547), .C1(new_n591), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n578), .A2(KEYINPUT29), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n572), .A2(new_n573), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n379), .B1(new_n563), .B2(new_n564), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n568), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT28), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT71), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT71), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n608), .A3(KEYINPUT28), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n603), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n601), .B1(new_n610), .B2(G902), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n568), .B1(new_n594), .B2(new_n581), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT29), .B1(new_n612), .B2(new_n579), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT70), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n566), .A2(new_n578), .A3(new_n572), .A4(new_n573), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n569), .B1(new_n604), .B2(new_n568), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT71), .ZN(new_n618));
  OAI211_X1 g432(.A(KEYINPUT72), .B(new_n254), .C1(new_n618), .C2(new_n603), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n613), .A2(new_n615), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT70), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n611), .A2(new_n616), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n600), .B1(new_n622), .B2(G472), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n574), .A2(new_n579), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n589), .A2(new_n590), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n599), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n546), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT69), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n547), .B1(new_n591), .B2(new_n599), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT69), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n545), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n544), .B1(new_n623), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT77), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT77), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n635), .B(new_n544), .C1(new_n623), .C2(new_n632), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n508), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n626), .A2(new_n254), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  INV_X1    g454(.A(new_n544), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n628), .A2(new_n640), .A3(new_n631), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n506), .B2(new_n507), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT33), .B1(new_n307), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n319), .A2(new_n320), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n645), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n309), .B2(new_n310), .ZN(new_n648));
  OAI21_X1  g462(.A(G478), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n312), .A2(new_n254), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n311), .B2(new_n312), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n645), .B1(new_n319), .B2(new_n320), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n309), .A2(new_n310), .A3(new_n647), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n312), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n312), .B(new_n254), .C1(new_n319), .C2(new_n320), .ZN(new_n657));
  INV_X1    g471(.A(new_n651), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT95), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n241), .A2(new_n244), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n426), .B(new_n258), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n643), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT34), .B(G104), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND2_X1  g484(.A1(new_n426), .A2(new_n258), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n663), .A2(new_n324), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n643), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT97), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n522), .A2(new_n523), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n527), .A3(new_n680), .ZN(new_n681));
  OAI22_X1  g495(.A1(new_n524), .A2(new_n528), .B1(KEYINPUT36), .B2(new_n512), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n678), .B1(new_n683), .B2(new_n541), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT98), .A4(new_n542), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n538), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n628), .A2(new_n640), .A3(new_n631), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n427), .ZN(new_n688));
  INV_X1    g502(.A(new_n507), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT85), .B1(new_n499), .B2(new_n503), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n687), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  NAND2_X1  g507(.A1(new_n506), .A2(new_n507), .ZN(new_n694));
  INV_X1    g508(.A(new_n686), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n623), .B2(new_n632), .ZN(new_n696));
  INV_X1    g510(.A(new_n251), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n698), .B2(new_n256), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n673), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n694), .A2(new_n696), .A3(new_n426), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(new_n699), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n694), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n663), .A2(new_n323), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n686), .A2(new_n709), .A3(new_n327), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  INV_X1    g525(.A(new_n600), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n596), .A2(new_n598), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n579), .B2(new_n605), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n714), .B2(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n632), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n424), .A2(new_n425), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n717), .B(new_n718), .Z(new_n719));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n271), .ZN(G45));
  AND3_X1   g540(.A1(new_n661), .A2(new_n663), .A3(new_n700), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n694), .A2(new_n696), .A3(new_n426), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  OAI21_X1  g543(.A(new_n254), .B1(new_n480), .B2(new_n486), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n503), .A3(new_n487), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n633), .A2(new_n667), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND3_X1  g550(.A1(new_n426), .A2(new_n258), .A3(new_n673), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n633), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n633), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  INV_X1    g558(.A(new_n325), .ZN(new_n745));
  AOI211_X1 g559(.A(new_n695), .B(new_n745), .C1(new_n623), .C2(new_n632), .ZN(new_n746));
  INV_X1    g560(.A(new_n487), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n432), .B1(new_n467), .B2(new_n468), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT84), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n479), .A3(new_n469), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n428), .B1(new_n751), .B2(new_n254), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n503), .A4(new_n426), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n731), .A2(new_n426), .A3(new_n503), .A4(new_n487), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  XNOR2_X1  g574(.A(new_n709), .B(KEYINPUT105), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n671), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n607), .A2(new_n609), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n572), .A2(new_n573), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n578), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n599), .A2(new_n625), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n546), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n640), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n641), .A3(new_n733), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  NAND4_X1  g584(.A1(new_n727), .A2(new_n640), .A3(new_n686), .A4(new_n767), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT106), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n758), .A2(new_n777), .A3(new_n772), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NOR2_X1   g594(.A1(new_n629), .A2(KEYINPUT32), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n781), .A2(new_n600), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n622), .A2(G472), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n781), .B2(new_n600), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n497), .B1(new_n495), .B2(KEYINPUT107), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(KEYINPUT107), .B2(new_n495), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n487), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n424), .A2(new_n503), .A3(new_n326), .A4(new_n425), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n661), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n792), .A2(new_n245), .A3(new_n793), .A4(new_n699), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n789), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n786), .A2(new_n795), .A3(new_n641), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n786), .A2(new_n795), .A3(KEYINPUT110), .A4(new_n641), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n623), .A2(new_n632), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n790), .B1(new_n788), .B2(new_n487), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n641), .A3(new_n727), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT108), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n793), .B1(new_n802), .B2(KEYINPUT108), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n798), .B(new_n799), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  NAND3_X1  g620(.A1(new_n633), .A2(new_n702), .A3(new_n801), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n633), .A2(new_n809), .A3(new_n702), .A4(new_n801), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G134), .ZN(G36));
  NAND2_X1  g626(.A1(new_n491), .A2(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n493), .A2(new_n494), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n816), .A3(G469), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT112), .A4(G469), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n496), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(KEYINPUT46), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n487), .B1(new_n821), .B2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n503), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n628), .A2(new_n640), .A3(new_n631), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n245), .A2(new_n661), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT43), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n827), .A2(KEYINPUT43), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n686), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT44), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n424), .A2(new_n326), .A3(new_n425), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n825), .A2(new_n832), .A3(new_n705), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  INV_X1    g650(.A(KEYINPUT47), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n824), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(KEYINPUT47), .B(new_n503), .C1(new_n822), .C2(new_n823), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n727), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n800), .A2(new_n641), .A3(new_n841), .A4(new_n833), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G140), .ZN(G42));
  XOR2_X1   g658(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n777), .B1(new_n758), .B2(new_n772), .ZN(new_n847));
  AOI211_X1 g661(.A(KEYINPUT106), .B(new_n771), .C1(new_n755), .C2(new_n757), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n717), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n761), .A2(new_n327), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n686), .A2(new_n502), .A3(new_n699), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n716), .A3(new_n789), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n703), .A2(new_n728), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n846), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n701), .B1(new_n506), .B2(new_n507), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n841), .B1(new_n506), .B2(new_n507), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n426), .B(new_n696), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n779), .A2(new_n858), .A3(KEYINPUT52), .A4(new_n853), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n633), .B(KEYINPUT77), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n861), .A2(new_n508), .B1(new_n742), .B2(new_n740), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n792), .A2(new_n245), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n672), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n323), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n318), .A2(new_n322), .A3(KEYINPUT113), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n663), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT114), .B1(new_n671), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n426), .A3(new_n872), .A4(new_n258), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n643), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n759), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n734), .A2(new_n691), .A3(new_n769), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n772), .A2(new_n801), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n245), .A2(new_n868), .A3(new_n700), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n881));
  INV_X1    g695(.A(new_n833), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n245), .A2(new_n868), .A3(new_n700), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT115), .B1(new_n884), .B2(new_n833), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n689), .B2(new_n690), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n800), .A2(new_n686), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n810), .B2(new_n808), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n805), .A2(new_n862), .A3(new_n878), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n845), .B1(new_n860), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n862), .A2(new_n878), .A3(new_n890), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n855), .A2(new_n859), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT53), .A4(new_n805), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n786), .A2(new_n641), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n829), .A2(new_n697), .A3(new_n828), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n900), .A2(new_n732), .A3(new_n833), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT48), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n716), .A2(new_n544), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n733), .A2(new_n697), .A3(new_n882), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n904), .A2(KEYINPUT120), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT120), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n906), .B(new_n907), .C1(new_n665), .C2(new_n664), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n247), .B(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n768), .A2(new_n641), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n900), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(new_n758), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n903), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n907), .A3(new_n245), .A4(new_n792), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n901), .A2(new_n686), .A3(new_n768), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n733), .A2(new_n327), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT118), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n910), .A2(new_n900), .A3(new_n719), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n918), .A2(KEYINPUT50), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT50), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n753), .A2(new_n502), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n838), .A2(new_n839), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n910), .A2(new_n900), .A3(new_n833), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n916), .B(new_n922), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT51), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n922), .B1(KEYINPUT119), .B2(KEYINPUT51), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n926), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT119), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(new_n916), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n913), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n860), .A2(new_n891), .A3(KEYINPUT117), .A4(new_n845), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n860), .A2(new_n891), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(KEYINPUT53), .ZN(new_n939));
  INV_X1    g753(.A(new_n845), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n936), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n898), .B(new_n935), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n246), .A2(new_n255), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n661), .A2(new_n245), .A3(new_n503), .A4(new_n326), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n731), .A2(new_n487), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n947), .B(new_n719), .C1(KEYINPUT49), .C2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(KEYINPUT49), .B2(new_n948), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(new_n904), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G75));
  NOR2_X1   g766(.A1(new_n255), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n254), .B1(new_n892), .B2(new_n895), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(G210), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n387), .A2(new_n390), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT123), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n408), .B(KEYINPUT55), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n896), .B2(G902), .ZN(new_n963));
  AOI211_X1 g777(.A(KEYINPUT124), .B(new_n254), .C1(new_n892), .C2(new_n895), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n423), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT56), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n966), .B2(new_n968), .ZN(G51));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n819), .A3(new_n820), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n496), .B(KEYINPUT57), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n943), .B1(new_n892), .B2(new_n895), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n897), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n751), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n953), .B1(new_n970), .B2(new_n974), .ZN(G54));
  INV_X1    g789(.A(new_n895), .ZN(new_n976));
  AND4_X1   g790(.A1(new_n805), .A2(new_n862), .A3(new_n878), .A4(new_n890), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n940), .B1(new_n977), .B2(new_n894), .ZN(new_n978));
  OAI21_X1  g792(.A(G902), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n955), .A2(new_n962), .ZN(new_n981));
  AND2_X1   g795(.A1(KEYINPUT58), .A2(G475), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n235), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n954), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n235), .B1(new_n965), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G60));
  NOR2_X1   g800(.A1(new_n646), .A2(new_n648), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n651), .B(KEYINPUT59), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n897), .B2(new_n972), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n954), .ZN(new_n992));
  INV_X1    g806(.A(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT53), .B1(new_n977), .B2(new_n894), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n941), .B1(KEYINPUT117), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n936), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n943), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n993), .B1(new_n997), .B2(new_n897), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n992), .B1(new_n998), .B2(new_n988), .ZN(G63));
  XOR2_X1   g813(.A(new_n533), .B(KEYINPUT60), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n896), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n539), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n1003), .B(new_n954), .C1(new_n683), .C2(new_n1001), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n953), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(KEYINPUT61), .C1(new_n683), .C2(new_n1001), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(G66));
  AND3_X1   g823(.A1(new_n734), .A2(new_n691), .A3(new_n769), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n746), .A2(new_n758), .B1(new_n643), .B2(new_n874), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1010), .A2(new_n743), .A3(new_n637), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(G953), .ZN(new_n1015));
  INV_X1    g829(.A(new_n253), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n1016), .B2(new_n406), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1015), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n958), .B1(G898), .B2(new_n255), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(G69));
  NAND4_X1  g838(.A1(new_n825), .A2(new_n705), .A3(new_n899), .A4(new_n851), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n835), .A2(new_n1025), .A3(new_n811), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n779), .A2(new_n858), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1027), .B1(new_n840), .B2(new_n842), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1026), .A2(new_n805), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n255), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n581), .B1(KEYINPUT30), .B2(new_n587), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n212), .A2(new_n213), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(G900), .B2(G953), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(KEYINPUT127), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(KEYINPUT62), .B1(new_n725), .B2(new_n1027), .ZN(new_n1040));
  INV_X1    g854(.A(new_n861), .ZN(new_n1041));
  INV_X1    g855(.A(new_n706), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1042), .B(new_n882), .C1(new_n863), .C2(new_n869), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n843), .B(new_n835), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  AND2_X1   g859(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  OR3_X1    g860(.A1(new_n725), .A2(KEYINPUT62), .A3(new_n1027), .ZN(new_n1047));
  AOI21_X1  g861(.A(G953), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1033), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1037), .B(new_n1039), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1047), .A2(new_n1045), .A3(new_n1040), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1049), .B1(new_n1051), .B2(new_n255), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1038), .B1(new_n1052), .B2(new_n1036), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1050), .A2(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(new_n612), .A2(new_n578), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1046), .A2(new_n1014), .A3(new_n1047), .ZN(new_n1056));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XOR2_X1   g871(.A(new_n1057), .B(KEYINPUT63), .Z(new_n1058));
  AOI21_X1  g872(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(new_n1058), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1060), .B1(new_n1029), .B2(new_n1014), .ZN(new_n1061));
  OR2_X1    g875(.A1(new_n612), .A2(new_n578), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n954), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n713), .B1(new_n579), .B2(new_n612), .ZN(new_n1064));
  NOR3_X1   g878(.A1(new_n942), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1059), .A2(new_n1063), .A3(new_n1065), .ZN(G57));
endmodule


