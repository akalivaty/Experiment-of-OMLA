//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT67), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n219), .A2(new_n220), .B1(G50), .B2(G226), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G68), .A2(G238), .ZN(new_n223));
  OAI21_X1  g0023(.A(KEYINPUT67), .B1(new_n214), .B2(new_n218), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n205), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n212), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  INV_X1    g0036(.A(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n202), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  XNOR2_X1  g0053(.A(KEYINPUT69), .B(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT70), .B(G223), .Z(new_n262));
  OAI211_X1 g0062(.A(new_n255), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n257), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n266), .C1(G77), .C2(new_n260), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n265), .A2(new_n269), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n267), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT71), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n279), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n230), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT72), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n278), .A2(new_n280), .A3(new_n283), .A4(new_n230), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT8), .B(G58), .Z(new_n290));
  NOR2_X1   g0090(.A1(new_n257), .A2(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n290), .A2(new_n291), .B1(G150), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n204), .B2(new_n231), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n231), .A2(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G13), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n289), .A2(new_n294), .B1(new_n202), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n282), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT73), .B1(new_n282), .B2(new_n284), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n299), .A2(new_n300), .A3(new_n295), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n275), .B1(new_n276), .B2(new_n274), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT9), .B1(new_n298), .B2(new_n302), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n274), .A2(G179), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n274), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n303), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n260), .A2(new_n254), .A3(G232), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G107), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n261), .B1(new_n258), .B2(new_n259), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G238), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n316), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n266), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n273), .A2(new_n226), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n271), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT15), .B(G87), .Z(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n291), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT76), .ZN(new_n333));
  INV_X1    g0133(.A(new_n290), .ZN(new_n334));
  INV_X1    g0134(.A(new_n292), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(new_n231), .B2(new_n205), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n285), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n297), .A2(new_n205), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n285), .A2(new_n295), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n276), .B2(new_n328), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n309), .B(new_n314), .C1(new_n330), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n328), .A2(new_n312), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n325), .A2(new_n346), .A3(new_n271), .A4(new_n327), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n254), .A2(G226), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G232), .A2(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n260), .ZN(new_n353));
  AND2_X1   g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n265), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n273), .A2(KEYINPUT77), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n265), .A2(new_n358), .A3(new_n269), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(G238), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n271), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT13), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n319), .B1(new_n350), .B2(new_n351), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n266), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n271), .A4(new_n360), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n366), .A3(KEYINPUT78), .ZN(new_n367));
  INV_X1    g0167(.A(new_n361), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n365), .A4(new_n364), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(G169), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n362), .A2(new_n366), .A3(KEYINPUT79), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT79), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(new_n374), .A3(new_n365), .A4(new_n364), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G179), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n367), .A2(new_n378), .A3(G169), .A4(new_n370), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n339), .A2(G68), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n296), .B2(G68), .ZN(new_n383));
  INV_X1    g0183(.A(G68), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n297), .A2(KEYINPUT12), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT80), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT80), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(new_n388), .A3(new_n383), .A4(new_n385), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n384), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n202), .B2(new_n335), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n289), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT11), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT11), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n289), .A2(new_n394), .A3(new_n391), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n387), .A2(new_n389), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n349), .B1(new_n380), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n254), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G87), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n399), .A2(new_n319), .B1(new_n257), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n266), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n265), .A2(G232), .A3(new_n269), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n271), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G190), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n290), .A2(new_n296), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n301), .B2(new_n290), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(G200), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n260), .B2(G20), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n317), .A2(new_n318), .A3(new_n410), .A4(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT81), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(G68), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(G58), .B(G68), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n384), .B1(new_n411), .B2(new_n413), .ZN(new_n422));
  INV_X1    g0222(.A(new_n419), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n285), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n406), .A2(new_n408), .A3(new_n409), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n408), .A2(new_n425), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n402), .A2(G179), .A3(new_n403), .A4(new_n271), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n405), .B2(new_n312), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n398), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n376), .A2(G190), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n367), .A2(G200), .A3(new_n370), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n396), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G107), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n216), .A2(new_n439), .A3(KEYINPUT6), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT82), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT6), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G97), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n441), .B1(new_n440), .B2(new_n443), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n440), .A2(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n444), .A3(G107), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n231), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT7), .B1(new_n319), .B2(new_n231), .ZN(new_n452));
  OAI21_X1  g0252(.A(G107), .B1(new_n452), .B2(new_n415), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n292), .A2(G77), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n285), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n297), .A2(new_n216), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n268), .A2(G33), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n287), .A2(new_n296), .A3(new_n288), .A4(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(new_n457), .C1(new_n216), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n463));
  OAI21_X1  g0263(.A(G244), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n464), .B2(new_n319), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n260), .A2(new_n254), .A3(KEYINPUT4), .A4(G244), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n321), .A2(G250), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n266), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n268), .B(G45), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n265), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n268), .A2(G45), .ZN(new_n475));
  OR2_X1    g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NAND2_X1  g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G274), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT83), .B1(new_n474), .B2(new_n479), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n474), .A2(new_n479), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(new_n479), .A3(KEYINPUT83), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT84), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n346), .B(new_n470), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n470), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n312), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n460), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n470), .A2(G190), .A3(new_n486), .A4(new_n487), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n482), .B1(new_n480), .B2(new_n481), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(KEYINPUT84), .A3(new_n487), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n490), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G200), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n460), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G238), .B1(new_n462), .B2(new_n463), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G244), .A2(G1698), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n319), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n257), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n266), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n265), .A2(G250), .A3(new_n475), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n265), .A2(KEYINPUT86), .A3(G250), .A4(new_n475), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n475), .A2(new_n270), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n511), .A3(new_n276), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n511), .A3(new_n513), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(G200), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n331), .A2(new_n296), .ZN(new_n518));
  AOI21_X1  g0318(.A(G20), .B1(new_n258), .B2(new_n259), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G68), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n400), .A2(new_n216), .A3(new_n439), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(KEYINPUT19), .C1(G20), .C2(new_n354), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT19), .B1(new_n354), .B2(new_n231), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n518), .B1(new_n285), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n523), .B1(new_n519), .B2(G68), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n522), .A2(new_n529), .B1(new_n282), .B2(new_n284), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT87), .B1(new_n530), .B2(new_n518), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n299), .A2(new_n300), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(G87), .A3(new_n296), .A4(new_n458), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n517), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n459), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n331), .B1(new_n528), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n515), .A2(new_n312), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n506), .A2(new_n511), .A3(new_n346), .A4(new_n513), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n535), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n500), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n468), .B(new_n231), .C1(G33), .C2(new_n216), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n281), .B(new_n543), .C1(new_n231), .C2(G116), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n297), .A2(new_n504), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n296), .A2(G116), .A3(new_n458), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n285), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n462), .A2(new_n463), .ZN(new_n551));
  OAI221_X1 g0351(.A(new_n260), .B1(new_n237), .B2(new_n261), .C1(new_n551), .C2(new_n217), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n266), .C1(G303), .C2(new_n260), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n473), .A2(G270), .A3(new_n265), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n479), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(G169), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n296), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  AND2_X1   g0360(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n561));
  NOR2_X1   g0361(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n519), .A2(G87), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n231), .B(G87), .C1(new_n317), .C2(new_n318), .ZN(new_n565));
  OR2_X1    g0365(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n231), .A2(KEYINPUT23), .A3(G107), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n567), .A3(new_n572), .A4(KEYINPUT24), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n285), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n560), .B(new_n577), .C1(new_n459), .C2(new_n439), .ZN(new_n578));
  OAI21_X1  g0378(.A(G250), .B1(new_n462), .B2(new_n463), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n217), .A2(new_n261), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n319), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G294), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n257), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n266), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n473), .A2(G264), .A3(new_n265), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n479), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n312), .ZN(new_n588));
  INV_X1    g0388(.A(new_n586), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n580), .B1(new_n254), .B2(G250), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n590), .A2(new_n319), .B1(new_n257), .B2(new_n583), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n591), .B2(new_n266), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n346), .A3(new_n479), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n578), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n553), .A2(G179), .A3(new_n479), .A4(new_n554), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n550), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n550), .A2(KEYINPUT21), .A3(G169), .A4(new_n555), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n558), .A2(new_n594), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n550), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n555), .A2(G200), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n276), .C2(new_n555), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n592), .A2(new_n604), .A3(new_n276), .A4(new_n479), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n587), .A2(new_n498), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n585), .A2(new_n276), .A3(new_n479), .A4(new_n586), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT89), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT90), .B1(new_n609), .B2(new_n578), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n459), .A2(new_n439), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n577), .A2(new_n560), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n542), .A2(new_n600), .A3(new_n603), .A4(new_n617), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n344), .A2(new_n434), .A3(new_n438), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n314), .ZN(new_n620));
  INV_X1    g0420(.A(new_n433), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n398), .A2(new_n438), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n427), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT93), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(KEYINPUT93), .B1(new_n308), .B2(new_n307), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n344), .A2(new_n434), .A3(new_n438), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n456), .A2(new_n457), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n459), .A2(new_n216), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n494), .C1(new_n498), .C2(new_n497), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n536), .A2(G87), .B1(new_n528), .B2(new_n531), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n526), .A2(new_n527), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n530), .A2(KEYINPUT87), .A3(new_n518), .ZN(new_n634));
  INV_X1    g0434(.A(new_n331), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n633), .A2(new_n634), .B1(new_n459), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n540), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n632), .A2(new_n517), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n631), .A2(new_n638), .A3(new_n493), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n609), .A2(KEYINPUT90), .A3(new_n578), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT91), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n594), .B(KEYINPUT92), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n558), .A2(new_n598), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n597), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n499), .A2(new_n460), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n460), .A2(new_n489), .A3(new_n492), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n617), .A4(new_n638), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n643), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n537), .A2(new_n540), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n541), .B2(new_n493), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n638), .A2(new_n648), .A3(KEYINPUT26), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n627), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n626), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n558), .A2(new_n597), .A3(new_n598), .ZN(new_n661));
  INV_X1    g0461(.A(G13), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G20), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n268), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n601), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n661), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n603), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT94), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(KEYINPUT94), .A3(new_n603), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G330), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n617), .A2(new_n594), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n613), .B2(new_n670), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n594), .B2(new_n670), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n644), .A2(new_n669), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n661), .A2(new_n670), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n210), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n521), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n233), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n658), .A2(new_n670), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n658), .A2(KEYINPUT97), .A3(new_n670), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n649), .A2(new_n599), .A3(new_n617), .A4(new_n638), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n669), .B1(new_n657), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n490), .A2(new_n491), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n704), .B(new_n516), .C1(new_n596), .C2(KEYINPUT95), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n592), .B1(new_n595), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT96), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT96), .B(new_n710), .C1(new_n705), .C2(new_n707), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n497), .A2(G179), .A3(new_n516), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(new_n555), .A3(new_n587), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n669), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(KEYINPUT31), .C1(new_n618), .C2(new_n669), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n669), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n693), .B1(new_n722), .B2(G1), .ZN(G364));
  AND2_X1   g0523(.A1(new_n675), .A2(new_n676), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n663), .A2(G45), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n689), .A2(G1), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n677), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT98), .Z(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n230), .B1(G20), .B2(new_n312), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n249), .A2(G45), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n687), .A2(new_n260), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n234), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n736), .A2(new_n740), .B1(new_n504), .B2(new_n687), .ZN(new_n741));
  NAND3_X1  g0541(.A1(G355), .A2(new_n210), .A3(new_n260), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n735), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n231), .A2(new_n346), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n276), .A3(new_n498), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(G190), .A3(new_n498), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n205), .B1(new_n746), .B2(new_n248), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT99), .ZN(new_n748));
  INV_X1    g0548(.A(new_n744), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n276), .A3(new_n498), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n231), .B1(new_n752), .B2(G190), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n748), .B1(new_n202), .B2(new_n751), .C1(new_n216), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n498), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G20), .A3(new_n276), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n749), .A2(new_n498), .A3(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n260), .B1(new_n439), .B2(new_n756), .C1(new_n758), .C2(new_n384), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(G20), .A3(G190), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT100), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n400), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n752), .A2(G20), .A3(new_n276), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n754), .A2(new_n759), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  OR2_X1    g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  NAND2_X1  g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n758), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n767), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(new_n583), .B2(new_n753), .C1(new_n776), .C2(new_n745), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n750), .A2(G326), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n777), .A2(new_n778), .A3(new_n260), .ZN(new_n779));
  INV_X1    g0579(.A(new_n756), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n774), .B(new_n779), .C1(G283), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n764), .C1(new_n783), .C2(new_n746), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n771), .A2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n743), .B(new_n727), .C1(new_n785), .C2(new_n733), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n673), .A2(new_n732), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n729), .A2(new_n788), .ZN(G396));
  OAI22_X1  g0589(.A1(new_n343), .A2(new_n330), .B1(new_n342), .B2(new_n670), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n348), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n348), .A2(new_n669), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n658), .A2(new_n670), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n696), .A2(new_n698), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT104), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n791), .A2(new_n799), .A3(new_n793), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n796), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n720), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n727), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n794), .A2(new_n730), .ZN(new_n806));
  INV_X1    g0606(.A(new_n727), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n319), .B1(new_n766), .B2(new_n776), .C1(new_n758), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n753), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G97), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n756), .A2(new_n400), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n745), .A2(new_n504), .B1(new_n746), .B2(new_n583), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G303), .C2(new_n750), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n811), .B(new_n814), .C1(new_n439), .C2(new_n764), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT102), .Z(new_n816));
  INV_X1    g0616(.A(new_n746), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT103), .B(G143), .ZN(new_n818));
  INV_X1    g0618(.A(new_n745), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n758), .B2(new_n821), .C1(new_n822), .C2(new_n751), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n823), .A2(new_n824), .B1(G132), .B2(new_n767), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n248), .B2(new_n753), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n756), .A2(new_n384), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n764), .A2(new_n202), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n260), .B1(new_n823), .B2(new_n824), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n733), .B1(new_n816), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n733), .A2(new_n730), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n205), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n806), .A2(new_n807), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n805), .A2(new_n834), .ZN(G384));
  NAND2_X1  g0635(.A1(new_n796), .A2(new_n793), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n420), .A2(new_n289), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT16), .B1(new_n417), .B2(new_n419), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n295), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n533), .A2(new_n290), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n407), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n430), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n667), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n840), .B2(new_n844), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n847), .A3(new_n426), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT105), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT37), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n848), .B2(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n428), .A2(new_n846), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n431), .A2(new_n852), .A3(new_n426), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n847), .B1(new_n433), .B2(new_n427), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n837), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT105), .ZN(new_n859));
  INV_X1    g0659(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT37), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n433), .A2(new_n427), .ZN(new_n863));
  INV_X1    g0663(.A(new_n847), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n397), .A2(new_n669), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n437), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n380), .A2(new_n397), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n380), .A2(new_n397), .A3(new_n670), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n836), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n433), .A2(new_n846), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n854), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n852), .B1(new_n433), .B2(new_n427), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n837), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n866), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n872), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT106), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n875), .A2(new_n890), .A3(new_n877), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n879), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n699), .A2(new_n627), .A3(new_n702), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n626), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n862), .B2(new_n865), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n873), .A2(new_n794), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n716), .A3(new_n718), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n896), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n719), .A2(new_n884), .A3(KEYINPUT40), .A4(new_n900), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n902), .A2(new_n627), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(G330), .A3(new_n903), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n803), .A2(new_n627), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n904), .A2(new_n719), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n895), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n268), .B2(new_n663), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n447), .A2(new_n450), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n504), .B1(new_n910), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n232), .C1(KEYINPUT35), .C2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OAI21_X1  g0713(.A(G77), .B1(new_n248), .B2(new_n384), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n914), .A2(new_n233), .B1(G50), .B2(new_n384), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n662), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(G367));
  NAND2_X1  g0717(.A1(new_n679), .A2(new_n684), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n500), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT42), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n649), .B1(new_n630), .B2(new_n670), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n493), .B1(new_n921), .B2(new_n594), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n670), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n632), .A2(new_n670), .ZN(new_n924));
  MUX2_X1   g0724(.A(new_n653), .B(new_n638), .S(new_n924), .Z(new_n925));
  AOI22_X1  g0725(.A1(new_n920), .A2(new_n923), .B1(KEYINPUT43), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n682), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n921), .B1(new_n493), .B2(new_n670), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n928), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n685), .A2(new_n930), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT44), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n685), .A2(new_n930), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT45), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n682), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n929), .B1(new_n937), .B2(new_n935), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n918), .B1(new_n681), .B2(new_n684), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(new_n677), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n720), .A3(new_n703), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n722), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n688), .B(KEYINPUT41), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n726), .A2(G1), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n932), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n239), .A2(new_n738), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n735), .B(new_n952), .C1(new_n687), .C2(new_n331), .ZN(new_n953));
  INV_X1    g0753(.A(new_n764), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT107), .Z(new_n958));
  AOI22_X1  g0758(.A1(new_n757), .A2(G294), .B1(new_n819), .B2(G283), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n780), .A2(G97), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n782), .C2(new_n746), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G317), .B2(new_n767), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n319), .B1(new_n751), .B2(new_n776), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n955), .B2(new_n956), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n753), .A2(new_n439), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n753), .A2(new_n384), .ZN(new_n967));
  INV_X1    g0767(.A(G159), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n758), .A2(new_n968), .B1(new_n202), .B2(new_n745), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT108), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n970), .B2(new_n969), .C1(new_n205), .C2(new_n756), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n954), .A2(G58), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n767), .A2(G137), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n750), .A2(new_n818), .B1(new_n817), .B2(G150), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n973), .A2(new_n260), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n965), .A2(new_n966), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n953), .B1(new_n978), .B2(new_n733), .ZN(new_n979));
  INV_X1    g0779(.A(new_n732), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n979), .B(new_n807), .C1(new_n980), .C2(new_n925), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n951), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT109), .Z(G387));
  OAI221_X1 g0783(.A(new_n960), .B1(new_n202), .B2(new_n746), .C1(new_n821), .C2(new_n766), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n954), .A2(G77), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n810), .A2(new_n331), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n757), .A2(new_n290), .B1(new_n819), .B2(G68), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n985), .A2(new_n260), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n984), .B(new_n988), .C1(G159), .C2(new_n750), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT110), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n954), .A2(G294), .B1(G283), .B2(new_n810), .ZN(new_n991));
  INV_X1    g0791(.A(G317), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n745), .A2(new_n782), .B1(new_n746), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT111), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n776), .B2(new_n758), .C1(new_n783), .C2(new_n751), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT48), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n991), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n998), .A2(new_n999), .B1(new_n996), .B2(new_n995), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT49), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n260), .B1(new_n767), .B2(G326), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n504), .B2(new_n756), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n990), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(new_n733), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n681), .A2(new_n980), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n737), .B1(new_n244), .B2(new_n739), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n260), .A2(new_n210), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n690), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n290), .A2(new_n202), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  NAND2_X1  g0811(.A1(G68), .A2(G77), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1011), .A2(new_n739), .A3(new_n1012), .A4(new_n690), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n687), .A2(new_n439), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n735), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR4_X1   g0816(.A1(new_n1005), .A2(new_n727), .A3(new_n1006), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n950), .B2(new_n944), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n721), .A2(new_n943), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n688), .A3(new_n945), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(G393));
  OR2_X1    g0821(.A1(new_n930), .A2(new_n980), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n954), .A2(G68), .B1(new_n767), .B2(new_n818), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT113), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n757), .A2(G50), .B1(new_n819), .B2(new_n290), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n260), .B1(new_n205), .B2(new_n753), .C1(new_n1026), .C2(KEYINPUT114), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n812), .B(new_n1027), .C1(new_n1024), .C2(new_n1023), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n750), .A2(G150), .B1(new_n817), .B2(G159), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT51), .Z(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1025), .B(new_n1031), .C1(KEYINPUT114), .C2(new_n1026), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n260), .B1(new_n767), .B2(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n439), .B2(new_n756), .C1(new_n764), .C2(new_n808), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n750), .A2(G317), .B1(new_n817), .B2(G311), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G116), .B2(new_n810), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1035), .B(new_n1038), .C1(new_n583), .C2(new_n745), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G303), .B2(new_n757), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n733), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n734), .B1(new_n216), .B2(new_n210), .C1(new_n252), .C2(new_n738), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1022), .A2(new_n807), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n941), .A2(new_n945), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n946), .A2(new_n688), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT116), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n946), .A2(KEYINPUT116), .A3(new_n1045), .A4(new_n688), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n939), .A2(new_n940), .A3(new_n950), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(G390));
  NAND3_X1  g0852(.A1(new_n893), .A2(new_n626), .A3(new_n906), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n716), .A2(G330), .A3(new_n718), .A4(new_n795), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1055), .A2(new_n873), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n873), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n836), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1055), .A2(new_n873), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n792), .B1(new_n701), .B2(new_n791), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n801), .A2(G330), .A3(new_n716), .A4(new_n718), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n873), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1054), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT117), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n871), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n872), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n884), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n791), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n669), .B(new_n1071), .C1(new_n657), .C2(new_n700), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n871), .B1(new_n1072), .B2(new_n792), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1073), .A2(KEYINPUT117), .A3(new_n884), .A4(new_n872), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n669), .B(new_n794), .C1(new_n652), .C2(new_n657), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n874), .B1(new_n1076), .B2(new_n792), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(new_n872), .B1(new_n886), .B2(new_n888), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1057), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n886), .A2(new_n888), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n873), .B1(new_n796), .B2(new_n793), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n887), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(new_n1070), .A3(new_n1074), .A4(new_n1059), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1065), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1054), .A2(new_n1079), .A3(new_n1083), .A4(new_n1064), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n688), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1080), .A2(new_n730), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n832), .A2(new_n334), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT53), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n954), .B2(G150), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n821), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G132), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1094), .A2(new_n745), .B1(new_n1095), .B2(new_n746), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n260), .B1(new_n766), .B2(new_n1098), .C1(new_n756), .C2(new_n202), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT118), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G137), .B2(new_n757), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1097), .B(new_n1101), .C1(new_n968), .C2(new_n753), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G128), .B2(new_n750), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n745), .A2(new_n216), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n765), .A2(new_n260), .A3(new_n827), .A4(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n751), .A2(new_n808), .B1(new_n753), .B2(new_n205), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G107), .B2(new_n757), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n583), .C2(new_n766), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G116), .B2(new_n817), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n733), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1088), .A2(new_n807), .A3(new_n1089), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n950), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1084), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT119), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(KEYINPUT119), .B(new_n1111), .C1(new_n1084), .C2(new_n1112), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1087), .A2(new_n1115), .A3(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n1053), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1053), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(KEYINPUT106), .B(new_n876), .C1(new_n1081), .C2(new_n867), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n890), .B1(new_n875), .B2(new_n877), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n309), .A2(new_n314), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1127), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n309), .A2(new_n314), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n303), .A2(new_n846), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n303), .A3(new_n846), .A4(new_n1130), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n902), .A2(new_n1135), .A3(G330), .A4(new_n903), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n905), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1125), .A2(new_n889), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n892), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1118), .B1(new_n1122), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1054), .B1(new_n1084), .B2(new_n1120), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(KEYINPUT57), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n688), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n727), .B1(new_n1135), .B2(new_n730), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n780), .A2(G58), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n985), .A2(new_n264), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G97), .B2(new_n757), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n319), .B1(new_n766), .B2(new_n808), .C1(new_n746), .C2(new_n439), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n967), .B(new_n1151), .C1(G116), .C2(new_n750), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n635), .C2(new_n745), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT58), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n202), .B1(new_n317), .B2(G41), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT120), .Z(new_n1158));
  OAI22_X1  g0958(.A1(new_n758), .A2(new_n1095), .B1(new_n753), .B2(new_n821), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n764), .A2(new_n1094), .B1(new_n1160), .B2(new_n746), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(G137), .C2(new_n819), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1098), .B2(new_n751), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n780), .A2(G159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n257), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1167), .A2(new_n1168), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n733), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n832), .A2(new_n202), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1147), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1139), .A2(new_n1141), .A3(new_n950), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1146), .A2(new_n1173), .A3(new_n1174), .ZN(G375));
  AND3_X1   g0975(.A1(new_n1120), .A2(new_n1053), .A3(KEYINPUT122), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT122), .B1(new_n1120), .B2(new_n1053), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n948), .B(new_n1065), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1120), .A2(KEYINPUT123), .A3(new_n1112), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n260), .B1(new_n954), .B2(G97), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n750), .A2(G294), .B1(G77), .B2(new_n780), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n504), .C2(new_n758), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n746), .A2(new_n808), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n766), .A2(new_n782), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n986), .B1(new_n439), .B2(new_n745), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n746), .A2(new_n822), .B1(new_n753), .B2(new_n202), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G58), .B2(new_n780), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n821), .B2(new_n745), .C1(new_n968), .C2(new_n764), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n766), .A2(new_n1160), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n751), .A2(new_n1095), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n260), .B1(new_n758), .B2(new_n1094), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n733), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n807), .B(new_n1194), .C1(new_n874), .C2(new_n731), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n384), .B2(new_n832), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT123), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1064), .B2(new_n950), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1179), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1178), .A2(new_n1199), .ZN(G381));
  NOR3_X1   g1000(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1201));
  OR2_X1    g1001(.A1(G375), .A2(G378), .ZN(new_n1202));
  OR2_X1    g1002(.A1(G393), .A2(G396), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1202), .A2(G381), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(G407));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1202), .ZN(G409));
  INV_X1    g1006(.A(new_n982), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT109), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G390), .A2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1050), .A2(new_n1051), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G390), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n982), .C1(G390), .C2(new_n1209), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n668), .A2(G213), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1144), .A2(new_n948), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(G378), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(G375), .C2(G378), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1176), .A2(new_n1177), .B1(new_n1121), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1120), .A2(new_n1053), .A3(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT124), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(KEYINPUT124), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n688), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(G384), .A3(new_n1199), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1227), .B2(new_n1199), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1221), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT62), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1221), .A2(new_n1235), .A3(new_n1231), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1217), .A2(G2897), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT125), .Z(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1227), .A2(new_n1199), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1228), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1221), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1216), .B1(new_n1237), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1212), .A2(new_n1215), .A3(new_n1234), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT63), .B1(new_n1221), .B2(new_n1246), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1232), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1217), .B1(G375), .B2(G378), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1220), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1231), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1221), .A2(new_n1256), .A3(KEYINPUT63), .A4(new_n1231), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1251), .A2(KEYINPUT127), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT127), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1248), .B1(new_n1259), .B2(new_n1260), .ZN(G405));
  XNOR2_X1  g1061(.A(G375), .B(G378), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(new_n1231), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(new_n1216), .Z(G402));
endmodule


