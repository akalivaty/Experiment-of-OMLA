//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT18), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n211), .B2(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G29gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT90), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n210), .A3(new_n217), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT91), .B1(new_n223), .B2(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n225), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n224), .A2(new_n230), .B1(new_n233), .B2(new_n223), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n208), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n207), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n230), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n223), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n235), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n223), .B(new_n230), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n235), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n237), .A3(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n239), .A2(new_n247), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G1gat), .B(G29gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT0), .ZN(new_n253));
  XNOR2_X1  g052(.A(G57gat), .B(G85gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257));
  XOR2_X1   g056(.A(G113gat), .B(G120gat), .Z(new_n258));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n262), .A3(G120gat), .ZN(new_n263));
  INV_X1    g062(.A(G127gat), .ZN(new_n264));
  INV_X1    g063(.A(G134gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G127gat), .A2(G134gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n261), .B(new_n263), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(new_n261), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT70), .B(G134gat), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G127gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n267), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT71), .A4(new_n273), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G141gat), .B(G148gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G155gat), .ZN(new_n281));
  INV_X1    g080(.A(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(KEYINPUT2), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n284), .B(new_n283), .C1(new_n279), .C2(KEYINPUT2), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n278), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT4), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n289), .B(KEYINPUT3), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(new_n278), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n257), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n257), .A3(new_n301), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT39), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n256), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n278), .B(new_n290), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n301), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n306), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n307), .A2(KEYINPUT85), .A3(KEYINPUT40), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n304), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n306), .B1(new_n313), .B2(new_n302), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(new_n311), .A3(KEYINPUT40), .A4(new_n255), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n294), .A2(KEYINPUT78), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n278), .A2(new_n320), .A3(new_n293), .A4(new_n290), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n321), .A3(new_n292), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n297), .A2(new_n301), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n308), .B2(new_n301), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n297), .B1(new_n292), .B2(new_n294), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n255), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n311), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT40), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337));
  INV_X1    g136(.A(G211gat), .ZN(new_n338));
  INV_X1    g137(.A(G218gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n335), .B1(new_n340), .B2(new_n336), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT69), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n355), .A4(new_n350), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT69), .B1(new_n351), .B2(new_n352), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n356), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n353), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G169gat), .ZN(new_n363));
  INV_X1    g162(.A(G176gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n365), .A2(KEYINPUT26), .A3(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n362), .B(new_n367), .C1(KEYINPUT26), .C2(new_n366), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n360), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(KEYINPUT23), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n373), .B2(new_n366), .ZN(new_n374));
  NAND3_X1  g173(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(G183gat), .B2(G190gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n361), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(KEYINPUT25), .B(new_n371), .C1(new_n373), .C2(new_n366), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n361), .A2(KEYINPUT64), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n376), .B1(new_n386), .B2(KEYINPUT66), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n388), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n379), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n384), .A2(new_n388), .A3(new_n385), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n384), .B2(new_n385), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n393), .A2(new_n394), .A3(new_n376), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n395), .A2(KEYINPUT67), .A3(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n369), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n347), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n369), .B(new_n400), .C1(new_n392), .C2(new_n396), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT67), .B1(new_n395), .B2(new_n380), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n389), .ZN(new_n404));
  INV_X1    g203(.A(new_n380), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n391), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n406), .A3(new_n379), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n407), .B2(new_n369), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n347), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n399), .B1(new_n409), .B2(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n397), .A2(KEYINPUT76), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n346), .B1(new_n411), .B2(new_n401), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n345), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n398), .B(new_n346), .C1(new_n402), .C2(new_n408), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n407), .A2(new_n347), .A3(new_n369), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n344), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n415), .B2(new_n418), .ZN(new_n426));
  INV_X1    g225(.A(new_n399), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n412), .B2(new_n413), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n344), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n418), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n318), .A2(new_n334), .A3(new_n424), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n398), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n344), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n336), .A2(new_n340), .ZN(new_n442));
  INV_X1    g241(.A(new_n335), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n444), .B2(new_n341), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(KEYINPUT81), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n398), .B1(new_n342), .B2(new_n343), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n440), .B1(new_n450), .B2(new_n289), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n441), .B1(new_n445), .B2(KEYINPUT80), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n453), .B(KEYINPUT29), .C1(new_n444), .C2(new_n341), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n289), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n439), .B1(new_n455), .B2(new_n437), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n435), .B(G22gat), .C1(new_n451), .C2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT31), .B(G50gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n451), .A2(new_n456), .A3(G22gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g264(.A(G22gat), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT3), .B1(new_n447), .B2(new_n453), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n445), .A2(KEYINPUT80), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n290), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n437), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n438), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n289), .B1(new_n446), .B2(new_n449), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n439), .A3(new_n437), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n466), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n462), .B(new_n463), .C1(new_n465), .C2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n460), .B1(new_n464), .B2(new_n474), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n466), .A3(new_n473), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n435), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n461), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(KEYINPUT83), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n327), .A2(new_n255), .A3(new_n330), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n331), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT86), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n327), .A2(new_n330), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n256), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n327), .A2(new_n255), .A3(new_n330), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n488), .A2(KEYINPUT86), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n331), .A2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n494));
  AOI21_X1  g293(.A(new_n423), .B1(new_n419), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n345), .B1(new_n428), .B2(new_n429), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n416), .A2(new_n417), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n497), .B(KEYINPUT37), .C1(new_n345), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n493), .A2(new_n500), .A3(new_n432), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT37), .B1(new_n415), .B2(new_n418), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n496), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n434), .B(new_n482), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n397), .A2(new_n278), .ZN(new_n505));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n278), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n407), .A2(new_n508), .A3(new_n369), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT32), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT73), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G71gat), .ZN(new_n516));
  INV_X1    g315(.A(G99gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n510), .B(KEYINPUT32), .C1(new_n512), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n509), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n506), .ZN(new_n525));
  AOI211_X1 g324(.A(KEYINPUT34), .B(new_n507), .C1(new_n505), .C2(new_n509), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT75), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n519), .A3(new_n521), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(new_n528), .A3(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n537), .A3(new_n521), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n528), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT36), .A3(new_n531), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n485), .A2(KEYINPUT79), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n488), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n484), .A2(new_n543), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n433), .A2(new_n424), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(new_n482), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n504), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n534), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(new_n481), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n433), .A2(new_n424), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n475), .A3(new_n480), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n539), .B2(new_n528), .ZN(new_n556));
  AOI211_X1 g355(.A(KEYINPUT88), .B(new_n554), .C1(new_n546), .C2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n545), .A2(new_n544), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n552), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(KEYINPUT35), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n553), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n251), .B1(new_n548), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  AOI21_X1  g363(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT99), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G99gat), .B(G106gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n223), .A2(new_n231), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n231), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n220), .A2(new_n222), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G190gat), .B(G218gat), .Z(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n568), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n566), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n596));
  INV_X1    g395(.A(G71gat), .ZN(new_n597));
  INV_X1    g396(.A(G78gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(KEYINPUT94), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n600), .B1(new_n599), .B2(new_n594), .ZN(new_n604));
  INV_X1    g403(.A(G57gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G64gat), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n603), .B(new_n604), .C1(KEYINPUT94), .C2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n596), .B1(new_n595), .B2(new_n601), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT96), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n230), .B1(new_n609), .B2(new_n610), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT97), .ZN(new_n622));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n622), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n592), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G230gat), .ZN(new_n632));
  INV_X1    g431(.A(G233gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n577), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n576), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638));
  INV_X1    g437(.A(new_n609), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n576), .B(new_n636), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT101), .B1(new_n642), .B2(new_n609), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n578), .A2(new_n609), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n640), .A2(new_n641), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n578), .A2(new_n609), .A3(new_n641), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n634), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n634), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  OR2_X1    g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n647), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n634), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT102), .B1(new_n653), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n563), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n559), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(G1gat), .Z(G1324gat));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n229), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n663), .A2(new_n552), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n552), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n229), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT42), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n663), .B2(new_n542), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n549), .A2(G15gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n663), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n662), .A2(new_n481), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n628), .A2(new_n629), .ZN(new_n679));
  INV_X1    g478(.A(new_n592), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n680), .A3(new_n660), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n563), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n682), .A2(new_n211), .A3(new_n544), .A4(new_n545), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n504), .A2(new_n542), .A3(new_n547), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n562), .A2(KEYINPUT105), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(new_n553), .C1(new_n557), .C2(new_n561), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n693), .B2(new_n680), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n548), .A2(new_n562), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(KEYINPUT44), .A3(new_n592), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n679), .A2(new_n251), .A3(new_n660), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n559), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n686), .A2(new_n687), .A3(new_n700), .ZN(G1328gat));
  OAI21_X1  g500(.A(G36gat), .B1(new_n699), .B2(new_n552), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n682), .A2(new_n213), .A3(new_n669), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(new_n542), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G43gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n682), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n549), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n699), .A2(new_n707), .B1(G43gat), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n481), .A3(new_n696), .A4(new_n698), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n482), .A2(G50gat), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n682), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT106), .B1(new_n712), .B2(G50gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n713), .A2(new_n722), .A3(new_n716), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n713), .B2(new_n716), .ZN(new_n725));
  AOI211_X1 g524(.A(KEYINPUT107), .B(new_n715), .C1(new_n712), .C2(G50gat), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n725), .A2(new_n726), .B1(new_n720), .B2(new_n719), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n560), .A2(new_n558), .A3(KEYINPUT35), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n691), .B1(new_n732), .B2(new_n553), .ZN(new_n733));
  INV_X1    g532(.A(new_n692), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n548), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n631), .A2(new_n250), .A3(new_n659), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n559), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n605), .ZN(G1332gat));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n737), .B(new_n669), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n738), .A2(new_n552), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n741), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT108), .ZN(G1333gat));
  NAND3_X1  g545(.A1(new_n737), .A2(G71gat), .A3(new_n706), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT109), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n534), .B(KEYINPUT110), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n597), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT50), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n481), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n679), .A2(new_n250), .A3(new_n659), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n697), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n559), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n679), .A2(new_n250), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n592), .A4(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n690), .A2(new_n692), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n680), .B1(new_n765), .B2(new_n548), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n766), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n761), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n735), .A2(new_n592), .A3(new_n761), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n764), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n660), .A2(new_n573), .A3(new_n544), .A4(new_n545), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  NAND3_X1  g571(.A1(new_n660), .A2(new_n669), .A3(new_n574), .ZN(new_n773));
  AOI211_X1 g572(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n766), .C2(new_n761), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n769), .B2(new_n768), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n764), .A2(new_n767), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n694), .A2(new_n669), .A3(new_n696), .A4(new_n758), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n781), .C1(new_n770), .C2(new_n773), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n759), .B2(new_n542), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n660), .A2(new_n517), .A3(new_n534), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n770), .B2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n659), .A2(G106gat), .A3(new_n482), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n769), .A2(new_n768), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n778), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n694), .A2(new_n481), .A3(new_n696), .A4(new_n758), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n797), .B2(G106gat), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(KEYINPUT114), .C1(new_n770), .C2(new_n794), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n794), .B1(new_n777), .B2(new_n778), .ZN(new_n805));
  INV_X1    g604(.A(new_n798), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n243), .A2(new_n237), .A3(new_n207), .A4(new_n246), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n242), .A2(new_n235), .B1(new_n245), .B2(new_n244), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n206), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT117), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n592), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n810), .B2(new_n812), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n645), .A2(new_n634), .A3(new_n646), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n645), .A2(KEYINPUT115), .A3(new_n634), .A4(new_n646), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n654), .A3(KEYINPUT54), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n652), .B1(new_n647), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n656), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n656), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n826), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n828), .A2(new_n250), .A3(new_n826), .A4(new_n831), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n810), .A2(new_n812), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n657), .B2(new_n658), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n809), .B(new_n832), .C1(new_n836), .C2(new_n592), .ZN(new_n837));
  INV_X1    g636(.A(new_n679), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n592), .B1(new_n833), .B2(new_n835), .ZN(new_n839));
  INV_X1    g638(.A(new_n832), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n630), .A2(new_n251), .A3(new_n659), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n669), .A2(new_n559), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n481), .A3(new_n549), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n262), .B1(new_n847), .B2(new_n250), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT119), .Z(new_n849));
  INV_X1    g648(.A(new_n556), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n262), .A3(new_n250), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(G1340gat));
  AOI21_X1  g652(.A(G120gat), .B1(new_n851), .B2(new_n660), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n660), .A2(G120gat), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n847), .B2(new_n855), .ZN(G1341gat));
  AOI21_X1  g655(.A(new_n264), .B1(new_n847), .B2(new_n679), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n838), .A2(G127gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT120), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n680), .A2(new_n271), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT56), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n680), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n265), .B1(new_n864), .B2(new_n550), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n863), .A2(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(G141gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n542), .A2(new_n845), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n250), .A2(new_n656), .A3(new_n824), .A4(new_n831), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n592), .B1(new_n835), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n838), .B1(new_n840), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n482), .B1(new_n872), .B2(new_n843), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n482), .B1(new_n842), .B2(new_n843), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n874), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n867), .B1(new_n877), .B2(new_n250), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n876), .A2(new_n869), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n251), .A2(G141gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT58), .B1(new_n878), .B2(KEYINPUT121), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1344gat));
  INV_X1    g682(.A(G148gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n884), .A3(new_n660), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n876), .A2(new_n887), .A3(KEYINPUT57), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n876), .B2(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n660), .A3(new_n869), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n884), .C1(new_n877), .C2(new_n660), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n281), .A3(new_n679), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n877), .A2(new_n679), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n281), .ZN(G1346gat));
  NOR2_X1   g697(.A1(new_n706), .A2(new_n482), .ZN(new_n899));
  AOI21_X1  g698(.A(G162gat), .B1(new_n864), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n680), .A2(new_n282), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n877), .B2(new_n901), .ZN(G1347gat));
  NAND2_X1  g701(.A1(new_n669), .A2(new_n559), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n749), .A2(new_n903), .A3(new_n481), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n844), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n363), .A3(new_n251), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n844), .A2(new_n559), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT123), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n844), .A2(new_n909), .A3(new_n559), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n669), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n850), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n250), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n906), .B1(new_n913), .B2(new_n363), .ZN(G1348gat));
  NOR3_X1   g713(.A1(new_n905), .A2(new_n364), .A3(new_n659), .ZN(new_n915));
  AOI21_X1  g714(.A(G176gat), .B1(new_n912), .B2(new_n660), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1349gat));
  OAI21_X1  g718(.A(G183gat), .B1(new_n905), .B2(new_n838), .ZN(new_n920));
  INV_X1    g719(.A(new_n912), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n679), .A2(new_n349), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n905), .B2(new_n680), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n592), .A2(new_n350), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n921), .B2(new_n927), .ZN(G1351gat));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n669), .A3(new_n899), .A4(new_n910), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(KEYINPUT125), .B(G197gat), .Z(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n250), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n876), .A2(new_n887), .A3(KEYINPUT57), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n706), .A2(new_n903), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n874), .B(new_n482), .C1(new_n842), .C2(new_n843), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n933), .B(new_n934), .C1(new_n935), .C2(new_n889), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n251), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n937), .B2(new_n931), .ZN(G1352gat));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n891), .A2(KEYINPUT126), .A3(new_n660), .A4(new_n934), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n936), .B2(new_n659), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n940), .A2(new_n942), .A3(G204gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n659), .A2(G204gat), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n929), .A2(KEYINPUT62), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n929), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n939), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n940), .A2(new_n942), .A3(G204gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n950), .A2(KEYINPUT127), .A3(new_n947), .A4(new_n946), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n930), .A2(new_n338), .A3(new_n679), .ZN(new_n953));
  OAI21_X1  g752(.A(G211gat), .B1(new_n936), .B2(new_n838), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n936), .B2(new_n680), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n592), .A2(new_n339), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n929), .B2(new_n960), .ZN(G1355gat));
endmodule


