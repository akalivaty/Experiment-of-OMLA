//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n469), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n474), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n470), .A2(G2105), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n479), .B1(new_n480), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n471), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n474), .A2(new_n490), .A3(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n495), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n500), .A2(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G88), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n500), .A2(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT69), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n503), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT70), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n519), .A2(new_n520), .A3(new_n507), .A4(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(G166));
  XNOR2_X1  g097(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n524), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT6), .B(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G51), .A3(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(new_n536), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(G168));
  NAND3_X1  g116(.A1(new_n536), .A2(G52), .A3(G543), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(G90), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT5), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G64), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n503), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n545), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n536), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n538), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n512), .B2(G56), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n503), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  AND2_X1   g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  NOR2_X1   g141(.A1(KEYINPUT6), .A2(G651), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n536), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n500), .B2(new_n501), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n512), .A2(new_n536), .A3(G91), .ZN(new_n578));
  AND4_X1   g153(.A1(KEYINPUT74), .A2(new_n572), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(G65), .B1(new_n546), .B2(new_n547), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(new_n575), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n506), .B2(G91), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT74), .B1(new_n582), .B2(new_n572), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n579), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  INV_X1    g161(.A(G166), .ZN(G303));
  NAND2_X1  g162(.A1(new_n506), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n503), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n538), .A2(new_n594), .B1(new_n553), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n503), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n538), .A2(new_n601), .B1(new_n553), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n538), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n546), .A2(new_n547), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G321));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(G286), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G299), .B(KEYINPUT75), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G297));
  AOI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n618), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NAND2_X1  g207(.A1(new_n474), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n467), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n633), .B1(new_n634), .B2(new_n635), .C1(new_n636), .C2(new_n483), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT77), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n470), .A2(new_n468), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n649), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n674), .A2(new_n677), .A3(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT80), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G16), .A2(G22), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G166), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G1971), .Z(new_n694));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G6), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n597), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n698), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n696), .A2(new_n697), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n698), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n604), .B2(new_n698), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT82), .B(G1986), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT81), .ZN(new_n718));
  INV_X1    g293(.A(new_n483), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n474), .A2(G131), .ZN(new_n721));
  OR2_X1    g296(.A1(G95), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n716), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n710), .A2(new_n711), .A3(new_n715), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(KEYINPUT85), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n719), .A2(G129), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n716), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT90), .B2(new_n739), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(G160), .A2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n745), .B2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(KEYINPUT24), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n698), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n698), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT91), .Z(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n749), .B1(G1961), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n618), .B2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT86), .B(G1348), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n698), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n559), .B2(new_n698), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT87), .B(G1341), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n716), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n719), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n474), .A2(G140), .ZN(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(new_n716), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n758), .A2(new_n762), .A3(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n754), .A2(KEYINPUT92), .B1(KEYINPUT88), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n470), .A2(G127), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n467), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n782), .A2(new_n783), .B1(new_n474), .B2(G139), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n778), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n778), .B2(new_n784), .ZN(new_n787));
  OAI21_X1  g362(.A(G29), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G33), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(G29), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G2072), .ZN(new_n791));
  INV_X1    g366(.A(G1961), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n752), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G2072), .B2(new_n790), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n748), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n698), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n698), .B2(G21), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT30), .B(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(KEYINPUT31), .A2(G11), .ZN(new_n802));
  NAND2_X1  g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n801), .A2(new_n716), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n637), .B2(new_n716), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n795), .A2(new_n799), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n716), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n716), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT93), .B(G2078), .Z(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  NAND4_X1  g385(.A1(new_n774), .A2(new_n794), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G20), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT23), .ZN(new_n814));
  INV_X1    g389(.A(G299), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n698), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n818), .B1(new_n773), .B2(KEYINPUT88), .C1(new_n754), .C2(KEYINPUT92), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n716), .A2(G35), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G162), .B2(new_n716), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2090), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n811), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n732), .A2(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND2_X1  g402(.A1(new_n618), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n538), .A2(new_n830), .B1(new_n553), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n512), .A2(G67), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n503), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n558), .A2(new_n555), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G56), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(G651), .B1(new_n838), .B2(new_n556), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n506), .A2(G81), .B1(new_n509), .B2(G43), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n506), .A2(G93), .B1(new_n509), .B2(G55), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n834), .B1(new_n613), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G651), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n829), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n841), .A2(new_n844), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n851), .A2(new_n854), .ZN(G145));
  INV_X1    g430(.A(new_n784), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT89), .B1(new_n856), .B2(new_n777), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n785), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n857), .B2(new_n785), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n769), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n493), .A2(new_n495), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n492), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT97), .B1(new_n786), .B2(new_n787), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n770), .A3(new_n859), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n862), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n862), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n737), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n867), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n863), .B1(new_n489), .B2(new_n491), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n737), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n862), .A2(new_n865), .A3(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G130), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n467), .A2(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n483), .A2(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G142), .B2(new_n474), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n641), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n725), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n870), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n486), .B(G160), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n637), .B(KEYINPUT96), .Z(new_n887));
  XOR2_X1   g462(.A(new_n886), .B(new_n887), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n884), .B1(new_n870), .B2(new_n876), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n870), .A2(new_n876), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n896), .A2(KEYINPUT98), .A3(new_n883), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n885), .B1(new_n891), .B2(KEYINPUT98), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n852), .A2(new_n621), .ZN(new_n903));
  NAND2_X1  g478(.A1(G290), .A2(new_n597), .ZN(new_n904));
  NAND2_X1  g479(.A1(G305), .A2(new_n604), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n517), .A2(new_n521), .A3(G288), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G288), .B1(new_n517), .B2(new_n521), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G166), .A2(new_n704), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n911), .A2(new_n907), .A3(new_n904), .A4(new_n905), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n912), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n910), .B2(new_n912), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  MUX2_X1   g493(.A(KEYINPUT102), .B(new_n914), .S(new_n918), .Z(new_n919));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n579), .B2(new_n583), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT74), .ZN(new_n922));
  INV_X1    g497(.A(new_n572), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n577), .A2(new_n578), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n582), .A2(KEYINPUT74), .A3(new_n572), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(KEYINPUT100), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(new_n618), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(G299), .A2(KEYINPUT100), .A3(new_n617), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(KEYINPUT41), .A3(new_n929), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n847), .B(new_n628), .ZN(new_n936));
  MUX2_X1   g511(.A(new_n931), .B(new_n935), .S(new_n936), .Z(new_n937));
  XNOR2_X1  g512(.A(new_n919), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n903), .B1(new_n938), .B2(new_n621), .ZN(G295));
  OAI21_X1  g514(.A(new_n903), .B1(new_n938), .B2(new_n621), .ZN(G331));
  OAI22_X1  g515(.A1(new_n535), .A2(new_n540), .B1(new_n545), .B2(new_n550), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n506), .A2(G89), .B1(new_n509), .B2(G51), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n506), .A2(new_n543), .B1(new_n509), .B2(G52), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n526), .A2(new_n531), .B1(new_n512), .B2(new_n533), .ZN(new_n944));
  INV_X1    g519(.A(new_n550), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n836), .A2(new_n941), .A3(new_n845), .A4(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n846), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(KEYINPUT103), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n933), .A2(new_n934), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT104), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n955), .A3(new_n947), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n847), .A2(KEYINPUT105), .A3(new_n941), .A4(new_n946), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(new_n930), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n933), .A2(new_n952), .A3(new_n960), .A4(new_n934), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n954), .A2(new_n917), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n954), .A2(new_n959), .A3(new_n961), .ZN(new_n966));
  INV_X1    g541(.A(new_n917), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n962), .A2(new_n963), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n952), .A2(new_n930), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n958), .A2(new_n933), .A3(new_n934), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(KEYINPUT106), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n935), .A2(new_n975), .A3(new_n958), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n917), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n969), .B(new_n970), .C1(new_n978), .C2(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n971), .B2(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n966), .A2(new_n967), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(new_n965), .A3(new_n963), .A4(new_n962), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT107), .A2(new_n980), .A3(KEYINPUT44), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n970), .B1(new_n964), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT107), .B1(new_n985), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n979), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(new_n979), .C1(new_n983), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(G397));
  NAND2_X1  g566(.A1(new_n582), .A2(new_n572), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT57), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n498), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT117), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT68), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n863), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n495), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1002), .B2(new_n492), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n995), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n469), .A2(new_n477), .A3(G40), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n865), .A2(new_n1008), .A3(new_n996), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n872), .B2(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1007), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1956), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n469), .A2(new_n477), .A3(G40), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n865), .A2(new_n996), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n498), .A2(new_n996), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(KEYINPUT110), .A3(new_n1018), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1015), .B(new_n1019), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n994), .B1(new_n1013), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1007), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1009), .A2(new_n995), .A3(new_n1010), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1348), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1009), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2067), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n618), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(new_n1016), .A3(new_n998), .A4(new_n1005), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n817), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1014), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n993), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1025), .A2(new_n1038), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1025), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(KEYINPUT61), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT61), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1025), .B(new_n1038), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT121), .B(G1996), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1036), .A2(KEYINPUT122), .A3(new_n1047), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n1029), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n558), .B(new_n555), .C1(KEYINPUT123), .C2(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1054), .B(new_n1055), .C1(KEYINPUT123), .C2(KEYINPUT59), .ZN(new_n1059));
  NOR4_X1   g634(.A1(new_n1028), .A2(new_n1030), .A3(KEYINPUT60), .A4(new_n617), .ZN(new_n1060));
  OR3_X1    g635(.A1(new_n1028), .A2(new_n618), .A3(new_n1030), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1031), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(KEYINPUT60), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1039), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1029), .A2(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n596), .A2(KEYINPUT114), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  OAI221_X1 g643(.A(new_n1068), .B1(new_n553), .B2(new_n595), .C1(new_n594), .C2(new_n538), .ZN(new_n1069));
  INV_X1    g644(.A(new_n593), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G1981), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT113), .B(G1981), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n597), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1072), .A2(new_n1080), .A3(KEYINPUT49), .A4(new_n1074), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1066), .A2(new_n1076), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n704), .A2(G1976), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1029), .A2(G8), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1029), .A2(G8), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1082), .A2(KEYINPUT118), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1034), .A2(G2090), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1036), .A2(G1971), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G303), .A2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1091), .A2(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1036), .A2(G1971), .B1(new_n1102), .B2(G2090), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1104), .B2(new_n1099), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1103), .A2(KEYINPUT112), .A3(new_n1098), .A4(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G2078), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1036), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1016), .B1(new_n1022), .B2(new_n1018), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT45), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1113));
  OR4_X1    g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(G2078), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1102), .A2(new_n792), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(G171), .B(KEYINPUT54), .Z(new_n1117));
  AOI22_X1  g692(.A1(new_n1109), .A2(new_n1110), .B1(new_n792), .B2(new_n1102), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1110), .B(G2078), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1019), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1116), .A2(new_n1117), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1100), .A2(new_n1107), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n798), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1026), .A2(new_n743), .A3(new_n1027), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n1127), .B2(G286), .ZN(new_n1128));
  AOI21_X1  g703(.A(G168), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(G8), .C1(new_n1127), .C2(G286), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1130), .A2(new_n1124), .A3(new_n1132), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1123), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1065), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1133), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1130), .A2(new_n1124), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(KEYINPUT62), .A3(new_n1138), .ZN(new_n1139));
  AND4_X1   g714(.A1(G171), .A2(new_n1100), .A3(new_n1107), .A4(new_n1116), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1134), .B2(new_n1133), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(G168), .A2(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1127), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1104), .A2(new_n1099), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1089), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1107), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT120), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1100), .A2(new_n1107), .A3(new_n1149), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1151), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(new_n1107), .A3(new_n1158), .A4(new_n1150), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1154), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1107), .A2(new_n1089), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1082), .A2(new_n1084), .A3(new_n704), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1074), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1066), .B(KEYINPUT116), .Z(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1136), .A2(new_n1143), .A3(new_n1160), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1017), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1167), .A2(new_n1007), .A3(KEYINPUT45), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n769), .B(G2067), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT109), .Z(new_n1171));
  XNOR2_X1  g746(.A(new_n737), .B(G1996), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n725), .A2(new_n727), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n725), .A2(new_n727), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1168), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  NAND2_X1  g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1168), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1166), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1168), .ZN(new_n1183));
  OR3_X1    g758(.A1(new_n1183), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT46), .B1(new_n1183), .B2(G1996), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1169), .A2(new_n737), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1184), .A2(new_n1185), .B1(new_n1168), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT47), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n769), .A2(G2067), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1183), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1177), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1183), .A2(new_n1178), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT48), .Z(new_n1194));
  AOI211_X1 g769(.A(new_n1188), .B(new_n1191), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1182), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n1198));
  NOR4_X1   g772(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n891), .A2(new_n890), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n888), .A3(new_n885), .ZN(new_n1201));
  OAI21_X1  g775(.A(new_n963), .B1(new_n1201), .B2(new_n893), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1202), .B2(new_n899), .ZN(new_n1203));
  OAI21_X1  g777(.A(new_n969), .B1(new_n978), .B2(KEYINPUT43), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1198), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1206));
  NAND4_X1  g780(.A1(new_n901), .A2(KEYINPUT126), .A3(new_n1206), .A4(new_n1199), .ZN(new_n1207));
  AND2_X1   g781(.A1(new_n1205), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(G225));
endmodule


