

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XOR2_X1 U326 ( .A(KEYINPUT79), .B(n540), .Z(n562) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U328 ( .A(KEYINPUT45), .B(n365), .Z(n295) );
  XNOR2_X1 U329 ( .A(n336), .B(n294), .ZN(n337) );
  XNOR2_X1 U330 ( .A(n338), .B(n337), .ZN(n340) );
  NOR2_X1 U331 ( .A1(n544), .A2(n460), .ZN(n531) );
  INV_X1 U332 ( .A(G120GAT), .ZN(n454) );
  XOR2_X1 U333 ( .A(n548), .B(KEYINPUT28), .Z(n516) );
  XOR2_X1 U334 ( .A(n413), .B(n412), .Z(n509) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1341GAT) );
  XOR2_X1 U337 ( .A(G92GAT), .B(G85GAT), .Z(n297) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n339) );
  XOR2_X1 U340 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n299) );
  XNOR2_X1 U341 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U343 ( .A(n339), .B(n300), .Z(n302) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n432) );
  XOR2_X1 U345 ( .A(G148GAT), .B(G78GAT), .Z(n317) );
  XNOR2_X1 U346 ( .A(n432), .B(n317), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n309) );
  XOR2_X1 U348 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n304) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n305), .B(KEYINPUT73), .Z(n307) );
  XOR2_X1 U352 ( .A(G176GAT), .B(G64GAT), .Z(n422) );
  XOR2_X1 U353 ( .A(G57GAT), .B(KEYINPUT13), .Z(n352) );
  XNOR2_X1 U354 ( .A(n422), .B(n352), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n309), .B(n308), .Z(n458) );
  XOR2_X1 U357 ( .A(KEYINPUT41), .B(n458), .Z(n535) );
  XNOR2_X1 U358 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(KEYINPUT92), .ZN(n311) );
  XOR2_X1 U360 ( .A(n311), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(G155GAT), .ZN(n312) );
  XOR2_X1 U362 ( .A(n313), .B(n312), .Z(n391) );
  XOR2_X1 U363 ( .A(KEYINPUT95), .B(KEYINPUT90), .Z(n315) );
  XNOR2_X1 U364 ( .A(KEYINPUT91), .B(KEYINPUT94), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n316), .B(G106GAT), .Z(n319) );
  XNOR2_X1 U367 ( .A(G22GAT), .B(n317), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n391), .B(n320), .Z(n331) );
  XOR2_X1 U370 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n322) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U373 ( .A(n323), .B(KEYINPUT22), .Z(n329) );
  XOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT76), .Z(n325) );
  XNOR2_X1 U375 ( .A(G50GAT), .B(G218GAT), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n344) );
  XOR2_X1 U377 ( .A(G204GAT), .B(G211GAT), .Z(n327) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n414) );
  XNOR2_X1 U380 ( .A(n344), .B(n414), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n548) );
  INV_X1 U383 ( .A(KEYINPUT36), .ZN(n347) );
  XOR2_X1 U384 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n333) );
  XOR2_X1 U385 ( .A(G134GAT), .B(KEYINPUT77), .Z(n405) );
  XOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .Z(n415) );
  XNOR2_X1 U387 ( .A(n405), .B(n415), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U389 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U390 ( .A(KEYINPUT9), .B(KEYINPUT78), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT7), .Z(n342) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(n343), .Z(n379) );
  XNOR2_X1 U397 ( .A(n379), .B(n344), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n540) );
  XNOR2_X1 U399 ( .A(n347), .B(n562), .ZN(n586) );
  XOR2_X1 U400 ( .A(G155GAT), .B(G71GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(G8GAT), .B(G183GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U403 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n351) );
  XNOR2_X1 U404 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U406 ( .A(n352), .B(G78GAT), .Z(n354) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G127GAT), .Z(n431) );
  XNOR2_X1 U408 ( .A(n431), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n359), .B(KEYINPUT80), .Z(n362) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G1GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n360), .B(KEYINPUT71), .ZN(n371) );
  XNOR2_X1 U416 ( .A(n371), .B(KEYINPUT15), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n523) );
  INV_X1 U419 ( .A(n523), .ZN(n581) );
  NOR2_X1 U420 ( .A1(n586), .A2(n581), .ZN(n365) );
  NOR2_X1 U421 ( .A1(n458), .A2(n295), .ZN(n382) );
  XOR2_X1 U422 ( .A(G113GAT), .B(G15GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G141GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n368), .B(G50GAT), .Z(n370) );
  XOR2_X1 U426 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XNOR2_X1 U427 ( .A(n423), .B(G36GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U429 ( .A(n371), .B(KEYINPUT68), .Z(n373) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U433 ( .A(KEYINPUT30), .B(KEYINPUT72), .Z(n377) );
  XNOR2_X1 U434 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n521) );
  INV_X1 U438 ( .A(n521), .ZN(n570) );
  NAND2_X1 U439 ( .A1(n382), .A2(n570), .ZN(n388) );
  NAND2_X1 U440 ( .A1(n535), .A2(n521), .ZN(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT46), .B(n383), .ZN(n384) );
  NAND2_X1 U442 ( .A1(n384), .A2(n581), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n540), .A2(n385), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n386), .B(KEYINPUT47), .ZN(n387) );
  NAND2_X1 U445 ( .A1(n388), .A2(n387), .ZN(n390) );
  XOR2_X1 U446 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n544) );
  INV_X1 U448 ( .A(n391), .ZN(n413) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n393) );
  XNOR2_X1 U450 ( .A(KEYINPUT98), .B(KEYINPUT1), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n395) );
  XNOR2_X1 U453 ( .A(G1GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U455 ( .A(n397), .B(n396), .Z(n411) );
  XOR2_X1 U456 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n399) );
  XNOR2_X1 U457 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n435) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(n435), .Z(n401) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U462 ( .A(G148GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U463 ( .A(G120GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(n404), .B(G85GAT), .Z(n407) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(n405), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n419) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(G92GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U479 ( .A(G183GAT), .B(KEYINPUT86), .Z(n427) );
  XNOR2_X1 U480 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U482 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n428) );
  XOR2_X1 U483 ( .A(n429), .B(n428), .Z(n436) );
  XOR2_X1 U484 ( .A(n430), .B(n436), .Z(n543) );
  INV_X1 U485 ( .A(n543), .ZN(n512) );
  XNOR2_X1 U486 ( .A(n512), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U487 ( .A1(n509), .A2(n467), .ZN(n460) );
  XOR2_X1 U488 ( .A(G134GAT), .B(n431), .Z(n434) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U491 ( .A(n435), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U497 ( .A(KEYINPUT65), .B(KEYINPUT88), .Z(n444) );
  XNOR2_X1 U498 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n446) );
  XNOR2_X1 U501 ( .A(G190GAT), .B(G99GAT), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U503 ( .A(n448), .B(n447), .Z(n449) );
  XOR2_X1 U504 ( .A(n450), .B(n449), .Z(n463) );
  INV_X1 U505 ( .A(n463), .ZN(n550) );
  NAND2_X1 U506 ( .A1(n531), .A2(n550), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT111), .B(n451), .Z(n452) );
  NOR2_X1 U508 ( .A1(n516), .A2(n452), .ZN(n453) );
  XNOR2_X1 U509 ( .A(KEYINPUT112), .B(n453), .ZN(n527) );
  AND2_X1 U510 ( .A1(n535), .A2(n527), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n455) );
  INV_X1 U512 ( .A(n458), .ZN(n576) );
  NAND2_X1 U513 ( .A1(n521), .A2(n576), .ZN(n485) );
  NOR2_X1 U514 ( .A1(n562), .A2(n581), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT16), .ZN(n473) );
  NOR2_X1 U516 ( .A1(n516), .A2(n460), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT101), .B(n461), .Z(n462) );
  NAND2_X1 U518 ( .A1(n463), .A2(n462), .ZN(n472) );
  INV_X1 U519 ( .A(n509), .ZN(n547) );
  NAND2_X1 U520 ( .A1(n550), .A2(n512), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n548), .A2(n464), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n465), .Z(n469) );
  NOR2_X1 U523 ( .A1(n550), .A2(n548), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U525 ( .A1(n467), .A2(n568), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n547), .A2(n470), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n482) );
  NAND2_X1 U529 ( .A1(n473), .A2(n482), .ZN(n497) );
  NOR2_X1 U530 ( .A1(n485), .A2(n497), .ZN(n479) );
  NAND2_X1 U531 ( .A1(n479), .A2(n509), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n512), .A2(n479), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U537 ( .A1(n479), .A2(n550), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n479), .A2(n516), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT102), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NAND2_X1 U542 ( .A1(n581), .A2(n482), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n483), .A2(n586), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT37), .ZN(n508) );
  NOR2_X1 U545 ( .A1(n508), .A2(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n495) );
  NAND2_X1 U548 ( .A1(n495), .A2(n509), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n512), .A2(n495), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n493) );
  NAND2_X1 U555 ( .A1(n495), .A2(n550), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n495), .A2(n516), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n499) );
  NAND2_X1 U561 ( .A1(n570), .A2(n535), .ZN(n507) );
  NOR2_X1 U562 ( .A1(n507), .A2(n497), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n504), .A2(n509), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  XOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U567 ( .A1(n504), .A2(n512), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n550), .A2(n504), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n516), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n511) );
  NOR2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n509), .A2(n517), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1336GAT) );
  XOR2_X1 U578 ( .A(G92GAT), .B(KEYINPUT109), .Z(n514) );
  NAND2_X1 U579 ( .A1(n517), .A2(n512), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n550), .A2(n517), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n520), .Z(G1339GAT) );
  NAND2_X1 U587 ( .A1(n527), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n525) );
  NAND2_X1 U590 ( .A1(n527), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(G127GAT), .B(n526), .Z(G1342GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U594 ( .A1(n562), .A2(n527), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(G134GAT), .B(n530), .Z(G1343GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n568), .ZN(n539) );
  NOR2_X1 U598 ( .A1(n570), .A2(n539), .ZN(n532) );
  XOR2_X1 U599 ( .A(G141GAT), .B(n532), .Z(G1344GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n534) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n537) );
  INV_X1 U603 ( .A(n535), .ZN(n555) );
  NOR2_X1 U604 ( .A1(n555), .A2(n539), .ZN(n536) );
  XOR2_X1 U605 ( .A(n537), .B(n536), .Z(G1345GAT) );
  NOR2_X1 U606 ( .A1(n581), .A2(n539), .ZN(n538) );
  XOR2_X1 U607 ( .A(G155GAT), .B(n538), .Z(G1346GAT) );
  INV_X1 U608 ( .A(n539), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT54), .B(n545), .ZN(n546) );
  AND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n569) );
  NAND2_X1 U614 ( .A1(n548), .A2(n569), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT55), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n563) );
  NOR2_X1 U617 ( .A1(n570), .A2(n563), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n563), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n581), .A2(n563), .ZN(n561) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n561), .Z(G1350GAT) );
  INV_X1 U629 ( .A(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n585) );
  NOR2_X1 U635 ( .A1(n570), .A2(n585), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT60), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n585), .A2(n576), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n585), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n584) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

