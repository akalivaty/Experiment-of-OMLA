

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734;

  XNOR2_X1 U365 ( .A(n531), .B(n530), .ZN(n534) );
  INV_X1 U366 ( .A(G953), .ZN(n725) );
  XOR2_X1 U367 ( .A(n350), .B(n402), .Z(n343) );
  XOR2_X1 U368 ( .A(n453), .B(n452), .Z(n344) );
  NOR2_X1 U369 ( .A1(n526), .A2(n546), .ZN(n345) );
  NAND2_X2 U370 ( .A1(n667), .A2(n668), .ZN(n664) );
  INV_X2 U371 ( .A(n506), .ZN(n667) );
  XNOR2_X2 U372 ( .A(n411), .B(n410), .ZN(n497) );
  XNOR2_X2 U373 ( .A(n443), .B(n408), .ZN(n707) );
  XNOR2_X2 U374 ( .A(n365), .B(n364), .ZN(n443) );
  XOR2_X2 U375 ( .A(G104), .B(G107), .Z(n348) );
  OR2_X1 U376 ( .A1(KEYINPUT44), .A2(n732), .ZN(n567) );
  INV_X2 U377 ( .A(n554), .ZN(n584) );
  NOR2_X1 U378 ( .A1(n546), .A2(n545), .ZN(n548) );
  NOR2_X1 U379 ( .A1(n522), .A2(n495), .ZN(n643) );
  BUF_X1 U380 ( .A(n510), .Z(n577) );
  XNOR2_X1 U381 ( .A(n380), .B(G146), .ZN(n419) );
  NAND2_X1 U382 ( .A1(n369), .A2(n367), .ZN(n734) );
  AND2_X1 U383 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U384 ( .A(n562), .B(KEYINPUT33), .ZN(n684) );
  XNOR2_X1 U385 ( .A(n548), .B(n547), .ZN(n563) );
  XNOR2_X1 U386 ( .A(n519), .B(n518), .ZN(n653) );
  XNOR2_X1 U387 ( .A(n419), .B(n418), .ZN(n482) );
  XNOR2_X1 U388 ( .A(n374), .B(G143), .ZN(n469) );
  NAND2_X1 U389 ( .A1(n355), .A2(n540), .ZN(n721) );
  XNOR2_X2 U390 ( .A(n348), .B(n405), .ZN(n706) );
  NAND2_X1 U391 ( .A1(n393), .A2(n398), .ZN(n392) );
  NAND2_X1 U392 ( .A1(n345), .A2(n354), .ZN(n496) );
  AND2_X1 U393 ( .A1(n580), .A2(n352), .ZN(n354) );
  XNOR2_X1 U394 ( .A(n386), .B(KEYINPUT79), .ZN(n516) );
  NOR2_X1 U395 ( .A1(n383), .A2(n382), .ZN(n381) );
  OR2_X1 U396 ( .A1(n345), .A2(n385), .ZN(n384) );
  NAND2_X1 U397 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U398 ( .A1(n684), .A2(n346), .ZN(n378) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT15), .ZN(n594) );
  XNOR2_X1 U400 ( .A(n533), .B(n359), .ZN(n358) );
  AND2_X1 U401 ( .A1(n517), .A2(n516), .ZN(n360) );
  INV_X1 U402 ( .A(KEYINPUT46), .ZN(n359) );
  INV_X1 U403 ( .A(G125), .ZN(n380) );
  XNOR2_X1 U404 ( .A(n482), .B(n451), .ZN(n722) );
  XNOR2_X1 U405 ( .A(G116), .B(G107), .ZN(n463) );
  XNOR2_X1 U406 ( .A(n395), .B(n595), .ZN(n599) );
  INV_X1 U407 ( .A(KEYINPUT64), .ZN(n595) );
  NAND2_X1 U408 ( .A1(n392), .A2(n391), .ZN(n395) );
  NOR2_X1 U409 ( .A1(n377), .A2(n564), .ZN(n376) );
  NOR2_X1 U410 ( .A1(n574), .A2(n351), .ZN(n377) );
  NAND2_X1 U411 ( .A1(n561), .A2(n584), .ZN(n562) );
  XNOR2_X1 U412 ( .A(n414), .B(n413), .ZN(n546) );
  NAND2_X1 U413 ( .A1(n399), .A2(n459), .ZN(n526) );
  XNOR2_X1 U414 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U415 ( .A(n450), .B(KEYINPUT108), .ZN(n400) );
  XNOR2_X1 U416 ( .A(n475), .B(n474), .ZN(n522) );
  XNOR2_X1 U417 ( .A(n473), .B(KEYINPUT104), .ZN(n474) );
  INV_X1 U418 ( .A(KEYINPUT47), .ZN(n385) );
  INV_X1 U419 ( .A(n639), .ZN(n383) );
  NOR2_X1 U420 ( .A1(n657), .A2(n385), .ZN(n382) );
  XNOR2_X1 U421 ( .A(n361), .B(n441), .ZN(n723) );
  XNOR2_X1 U422 ( .A(n723), .B(G146), .ZN(n455) );
  XNOR2_X1 U423 ( .A(n407), .B(n406), .ZN(n442) );
  XNOR2_X1 U424 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n407) );
  XNOR2_X1 U425 ( .A(G116), .B(G113), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n366), .B(KEYINPUT3), .ZN(n365) );
  INV_X1 U427 ( .A(G119), .ZN(n366) );
  INV_X1 U428 ( .A(n594), .ZN(n394) );
  XNOR2_X1 U429 ( .A(n440), .B(KEYINPUT69), .ZN(n499) );
  INV_X1 U430 ( .A(KEYINPUT28), .ZN(n450) );
  NAND2_X1 U431 ( .A1(n499), .A2(n577), .ZN(n401) );
  XNOR2_X1 U432 ( .A(n507), .B(KEYINPUT1), .ZN(n554) );
  XNOR2_X1 U433 ( .A(n357), .B(n356), .ZN(n355) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n356) );
  XNOR2_X1 U435 ( .A(KEYINPUT73), .B(G110), .ZN(n405) );
  XNOR2_X1 U436 ( .A(n421), .B(n420), .ZN(n422) );
  INV_X1 U437 ( .A(KEYINPUT24), .ZN(n420) );
  XNOR2_X1 U438 ( .A(G119), .B(G110), .ZN(n421) );
  INV_X1 U439 ( .A(KEYINPUT10), .ZN(n418) );
  XNOR2_X1 U440 ( .A(n706), .B(n442), .ZN(n453) );
  XNOR2_X1 U441 ( .A(KEYINPUT16), .B(G122), .ZN(n408) );
  XNOR2_X1 U442 ( .A(n469), .B(KEYINPUT4), .ZN(n361) );
  BUF_X1 U443 ( .A(n554), .Z(n665) );
  NAND2_X1 U444 ( .A1(n587), .A2(KEYINPUT32), .ZN(n370) );
  NAND2_X1 U445 ( .A1(n372), .A2(KEYINPUT32), .ZN(n371) );
  NOR2_X1 U446 ( .A1(n514), .A2(n513), .ZN(n529) );
  XNOR2_X1 U447 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U448 ( .A(n389), .B(n387), .ZN(n624) );
  XNOR2_X1 U449 ( .A(n388), .B(n361), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n453), .B(n707), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n404), .B(n343), .ZN(n388) );
  AND2_X1 U452 ( .A1(n390), .A2(n396), .ZN(n689) );
  XNOR2_X1 U453 ( .A(n532), .B(KEYINPUT40), .ZN(n614) );
  NOR2_X1 U454 ( .A1(n379), .A2(n375), .ZN(n565) );
  NAND2_X1 U455 ( .A1(n378), .A2(n376), .ZN(n375) );
  XNOR2_X1 U456 ( .A(n570), .B(KEYINPUT94), .ZN(n571) );
  INV_X1 U457 ( .A(KEYINPUT31), .ZN(n570) );
  INV_X1 U458 ( .A(KEYINPUT93), .ZN(n575) );
  XNOR2_X1 U459 ( .A(n610), .B(n353), .ZN(n363) );
  AND2_X1 U460 ( .A1(n574), .A2(n351), .ZN(n346) );
  NOR2_X1 U461 ( .A1(n503), .A2(n665), .ZN(n347) );
  INV_X1 U462 ( .A(n498), .ZN(n519) );
  XOR2_X1 U463 ( .A(n448), .B(n447), .Z(n349) );
  XOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n350) );
  XNOR2_X1 U465 ( .A(KEYINPUT34), .B(KEYINPUT75), .ZN(n351) );
  XOR2_X1 U466 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n352) );
  XOR2_X1 U467 ( .A(n609), .B(KEYINPUT62), .Z(n353) );
  INV_X1 U468 ( .A(KEYINPUT2), .ZN(n396) );
  NAND2_X1 U469 ( .A1(n360), .A2(n358), .ZN(n357) );
  XNOR2_X1 U470 ( .A(n362), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U471 ( .A1(n363), .A2(n611), .ZN(n362) );
  NAND2_X1 U472 ( .A1(n368), .A2(n373), .ZN(n367) );
  NOR2_X1 U473 ( .A1(n587), .A2(KEYINPUT32), .ZN(n368) );
  INV_X1 U474 ( .A(n373), .ZN(n372) );
  NOR2_X1 U475 ( .A1(n587), .A2(n667), .ZN(n556) );
  AND2_X1 U476 ( .A1(n553), .A2(n506), .ZN(n373) );
  NAND2_X1 U477 ( .A1(n734), .A2(n636), .ZN(n560) );
  XNOR2_X2 U478 ( .A(G128), .B(KEYINPUT77), .ZN(n374) );
  NOR2_X1 U479 ( .A1(n684), .A2(n351), .ZN(n379) );
  XNOR2_X2 U480 ( .A(n510), .B(KEYINPUT6), .ZN(n582) );
  NOR2_X2 U481 ( .A1(n664), .A2(n507), .ZN(n573) );
  NAND2_X1 U482 ( .A1(n384), .A2(n381), .ZN(n386) );
  NAND2_X1 U483 ( .A1(n398), .A2(n397), .ZN(n390) );
  NAND2_X1 U484 ( .A1(n394), .A2(KEYINPUT2), .ZN(n391) );
  NOR2_X1 U485 ( .A1(n711), .A2(n594), .ZN(n393) );
  INV_X1 U486 ( .A(n711), .ZN(n397) );
  INV_X1 U487 ( .A(n721), .ZN(n398) );
  XNOR2_X2 U488 ( .A(n552), .B(KEYINPUT22), .ZN(n587) );
  BUF_X1 U489 ( .A(n697), .Z(n701) );
  XNOR2_X1 U490 ( .A(n558), .B(KEYINPUT85), .ZN(n559) );
  XNOR2_X1 U491 ( .A(n419), .B(n403), .ZN(n404) );
  INV_X1 U492 ( .A(KEYINPUT9), .ZN(n462) );
  INV_X1 U493 ( .A(G478), .ZN(n473) );
  XNOR2_X1 U494 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U495 ( .A(n722), .B(n422), .ZN(n427) );
  INV_X1 U496 ( .A(KEYINPUT42), .ZN(n527) );
  XNOR2_X1 U497 ( .A(n572), .B(n571), .ZN(n646) );
  XNOR2_X1 U498 ( .A(n528), .B(n527), .ZN(n733) );
  XNOR2_X1 U499 ( .A(KEYINPUT88), .B(KEYINPUT74), .ZN(n402) );
  NAND2_X1 U500 ( .A1(G224), .A2(n725), .ZN(n403) );
  INV_X1 U501 ( .A(G101), .ZN(n406) );
  NAND2_X1 U502 ( .A1(n624), .A2(n594), .ZN(n411) );
  INV_X1 U503 ( .A(G902), .ZN(n490) );
  INV_X1 U504 ( .A(G237), .ZN(n409) );
  NAND2_X1 U505 ( .A1(n490), .A2(n409), .ZN(n412) );
  AND2_X1 U506 ( .A1(n412), .A2(G210), .ZN(n410) );
  NAND2_X1 U507 ( .A1(n412), .A2(G214), .ZN(n652) );
  NAND2_X1 U508 ( .A1(n497), .A2(n652), .ZN(n414) );
  XNOR2_X1 U509 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n413) );
  XOR2_X1 U510 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n417) );
  NAND2_X1 U511 ( .A1(G234), .A2(n594), .ZN(n415) );
  XNOR2_X1 U512 ( .A(KEYINPUT20), .B(n415), .ZN(n428) );
  NAND2_X1 U513 ( .A1(G221), .A2(n428), .ZN(n416) );
  XNOR2_X1 U514 ( .A(n417), .B(n416), .ZN(n668) );
  XNOR2_X1 U515 ( .A(G137), .B(G140), .ZN(n451) );
  XOR2_X1 U516 ( .A(G128), .B(KEYINPUT23), .Z(n425) );
  NAND2_X1 U517 ( .A1(G234), .A2(n725), .ZN(n423) );
  XOR2_X1 U518 ( .A(KEYINPUT8), .B(n423), .Z(n467) );
  NAND2_X1 U519 ( .A1(G221), .A2(n467), .ZN(n424) );
  XNOR2_X1 U520 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U521 ( .A(n427), .B(n426), .ZN(n702) );
  NOR2_X1 U522 ( .A1(G902), .A2(n702), .ZN(n433) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n430) );
  NAND2_X1 U524 ( .A1(n428), .A2(G217), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U526 ( .A(KEYINPUT90), .B(n431), .ZN(n432) );
  XNOR2_X1 U527 ( .A(n433), .B(n432), .ZN(n505) );
  XOR2_X1 U528 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n435) );
  NAND2_X1 U529 ( .A1(G234), .A2(G237), .ZN(n434) );
  XNOR2_X1 U530 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U531 ( .A1(G952), .A2(n436), .ZN(n683) );
  NOR2_X1 U532 ( .A1(n683), .A2(G953), .ZN(n544) );
  NAND2_X1 U533 ( .A1(G902), .A2(n436), .ZN(n542) );
  OR2_X1 U534 ( .A1(n725), .A2(n542), .ZN(n437) );
  NOR2_X1 U535 ( .A1(n437), .A2(G900), .ZN(n438) );
  NOR2_X1 U536 ( .A1(n544), .A2(n438), .ZN(n508) );
  NOR2_X1 U537 ( .A1(n505), .A2(n508), .ZN(n439) );
  NAND2_X1 U538 ( .A1(n668), .A2(n439), .ZN(n440) );
  INV_X1 U539 ( .A(G134), .ZN(n612) );
  XNOR2_X1 U540 ( .A(n612), .B(G131), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n443), .B(n442), .ZN(n448) );
  NOR2_X1 U542 ( .A1(G953), .A2(G237), .ZN(n478) );
  NAND2_X1 U543 ( .A1(n478), .A2(G210), .ZN(n444) );
  XNOR2_X1 U544 ( .A(n444), .B(KEYINPUT72), .ZN(n446) );
  XNOR2_X1 U545 ( .A(KEYINPUT5), .B(G137), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U547 ( .A(n455), .B(n349), .ZN(n609) );
  OR2_X2 U548 ( .A1(n609), .A2(G902), .ZN(n449) );
  XNOR2_X2 U549 ( .A(n449), .B(G472), .ZN(n510) );
  INV_X1 U550 ( .A(n451), .ZN(n452) );
  NAND2_X1 U551 ( .A1(G227), .A2(n725), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n344), .B(n454), .ZN(n456) );
  XNOR2_X1 U553 ( .A(n456), .B(n455), .ZN(n602) );
  NAND2_X1 U554 ( .A1(n602), .A2(n490), .ZN(n458) );
  XOR2_X1 U555 ( .A(KEYINPUT70), .B(G469), .Z(n457) );
  XNOR2_X2 U556 ( .A(n458), .B(n457), .ZN(n507) );
  XNOR2_X1 U557 ( .A(n507), .B(KEYINPUT107), .ZN(n459) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n461) );
  XNOR2_X1 U559 ( .A(G122), .B(KEYINPUT103), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n461), .B(n460), .ZN(n465) );
  XOR2_X1 U561 ( .A(n466), .B(KEYINPUT101), .Z(n472) );
  NAND2_X1 U562 ( .A1(n467), .A2(G217), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n468), .B(G134), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n698) );
  NOR2_X1 U566 ( .A1(G902), .A2(n698), .ZN(n475) );
  XOR2_X1 U567 ( .A(KEYINPUT98), .B(G140), .Z(n477) );
  XNOR2_X1 U568 ( .A(G143), .B(G122), .ZN(n476) );
  XNOR2_X1 U569 ( .A(n477), .B(n476), .ZN(n480) );
  NAND2_X1 U570 ( .A1(n478), .A2(G214), .ZN(n479) );
  XNOR2_X1 U571 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U572 ( .A(n482), .B(n481), .ZN(n489) );
  XOR2_X1 U573 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n484) );
  XNOR2_X1 U574 ( .A(KEYINPUT97), .B(KEYINPUT12), .ZN(n483) );
  XNOR2_X1 U575 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U576 ( .A(n485), .B(G104), .Z(n487) );
  XNOR2_X1 U577 ( .A(G113), .B(G131), .ZN(n486) );
  XNOR2_X1 U578 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n489), .B(n488), .ZN(n616) );
  NAND2_X1 U580 ( .A1(n616), .A2(n490), .ZN(n494) );
  XOR2_X1 U581 ( .A(KEYINPUT100), .B(KEYINPUT13), .Z(n492) );
  XNOR2_X1 U582 ( .A(KEYINPUT99), .B(G475), .ZN(n491) );
  XOR2_X1 U583 ( .A(n492), .B(n491), .Z(n493) );
  XNOR2_X1 U584 ( .A(n494), .B(n493), .ZN(n521) );
  INV_X1 U585 ( .A(n521), .ZN(n495) );
  AND2_X1 U586 ( .A1(n522), .A2(n495), .ZN(n645) );
  OR2_X1 U587 ( .A1(n643), .A2(n645), .ZN(n657) );
  XNOR2_X1 U588 ( .A(KEYINPUT80), .B(n657), .ZN(n580) );
  XNOR2_X1 U589 ( .A(n496), .B(KEYINPUT71), .ZN(n504) );
  INV_X1 U590 ( .A(n497), .ZN(n498) );
  NAND2_X1 U591 ( .A1(n643), .A2(n499), .ZN(n500) );
  NOR2_X1 U592 ( .A1(n582), .A2(n500), .ZN(n501) );
  AND2_X1 U593 ( .A1(n501), .A2(n652), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n519), .A2(n537), .ZN(n502) );
  XNOR2_X1 U595 ( .A(n502), .B(KEYINPUT36), .ZN(n503) );
  NOR2_X1 U596 ( .A1(n504), .A2(n347), .ZN(n517) );
  INV_X1 U597 ( .A(n505), .ZN(n506) );
  INV_X1 U598 ( .A(n508), .ZN(n509) );
  NAND2_X1 U599 ( .A1(n573), .A2(n509), .ZN(n514) );
  NAND2_X1 U600 ( .A1(n510), .A2(n652), .ZN(n512) );
  XNOR2_X1 U601 ( .A(KEYINPUT106), .B(KEYINPUT30), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U603 ( .A1(n522), .A2(n521), .ZN(n564) );
  NOR2_X1 U604 ( .A1(n564), .A2(n498), .ZN(n515) );
  NAND2_X1 U605 ( .A1(n529), .A2(n515), .ZN(n639) );
  XOR2_X1 U606 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n525) );
  INV_X1 U607 ( .A(KEYINPUT38), .ZN(n518) );
  NAND2_X1 U608 ( .A1(n652), .A2(n653), .ZN(n520) );
  XNOR2_X2 U609 ( .A(n520), .B(KEYINPUT109), .ZN(n658) );
  NOR2_X1 U610 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n523), .B(KEYINPUT105), .ZN(n655) );
  INV_X1 U612 ( .A(n655), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n658), .A2(n550), .ZN(n524) );
  XNOR2_X1 U614 ( .A(n525), .B(n524), .ZN(n686) );
  NOR2_X1 U615 ( .A1(n686), .A2(n526), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n529), .A2(n653), .ZN(n531) );
  XOR2_X1 U617 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n530) );
  NAND2_X1 U618 ( .A1(n534), .A2(n643), .ZN(n532) );
  NAND2_X1 U619 ( .A1(n733), .A2(n614), .ZN(n533) );
  INV_X1 U620 ( .A(n534), .ZN(n536) );
  INV_X1 U621 ( .A(n645), .ZN(n535) );
  NOR2_X1 U622 ( .A1(n536), .A2(n535), .ZN(n613) );
  NAND2_X1 U623 ( .A1(n665), .A2(n537), .ZN(n538) );
  XNOR2_X1 U624 ( .A(n538), .B(KEYINPUT43), .ZN(n539) );
  AND2_X1 U625 ( .A1(n539), .A2(n498), .ZN(n651) );
  NOR2_X1 U626 ( .A1(n613), .A2(n651), .ZN(n540) );
  XOR2_X1 U627 ( .A(KEYINPUT76), .B(n582), .Z(n541) );
  NOR2_X1 U628 ( .A1(n665), .A2(n541), .ZN(n553) );
  OR2_X1 U629 ( .A1(n725), .A2(G898), .ZN(n710) );
  NOR2_X1 U630 ( .A1(n710), .A2(n542), .ZN(n543) );
  NOR2_X1 U631 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U632 ( .A(KEYINPUT86), .B(KEYINPUT0), .Z(n547) );
  INV_X1 U633 ( .A(n668), .ZN(n549) );
  NOR2_X1 U634 ( .A1(n563), .A2(n549), .ZN(n551) );
  NAND2_X1 U635 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U636 ( .A1(n584), .A2(n577), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n556), .A2(n555), .ZN(n636) );
  INV_X1 U638 ( .A(KEYINPUT44), .ZN(n557) );
  NAND2_X1 U639 ( .A1(n557), .A2(KEYINPUT84), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n560), .B(n559), .ZN(n566) );
  NOR2_X1 U641 ( .A1(n582), .A2(n664), .ZN(n561) );
  INV_X1 U642 ( .A(n563), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n565), .B(KEYINPUT35), .ZN(n732) );
  NAND2_X1 U644 ( .A1(n566), .A2(n732), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n591) );
  INV_X1 U646 ( .A(n577), .ZN(n672) );
  NOR2_X1 U647 ( .A1(n664), .A2(n672), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n584), .A2(n569), .ZN(n674) );
  NOR2_X1 U649 ( .A1(n563), .A2(n674), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(n575), .ZN(n578) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n632) );
  NOR2_X1 U653 ( .A1(n646), .A2(n632), .ZN(n579) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT95), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n589) );
  INV_X1 U656 ( .A(n582), .ZN(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n667), .A2(n585), .ZN(n586) );
  NOR2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n629) );
  INV_X1 U660 ( .A(n629), .ZN(n588) );
  AND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U662 ( .A(KEYINPUT45), .ZN(n592) );
  XNOR2_X2 U663 ( .A(n593), .B(n592), .ZN(n711) );
  INV_X1 U664 ( .A(n721), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n596), .A2(KEYINPUT2), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n597), .B(KEYINPUT82), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n598), .A2(n711), .ZN(n690) );
  NOR2_X2 U668 ( .A1(n599), .A2(n690), .ZN(n697) );
  NAND2_X1 U669 ( .A1(n697), .A2(G469), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT57), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U674 ( .A(G952), .ZN(n605) );
  AND2_X1 U675 ( .A1(n605), .A2(G953), .ZN(n705) );
  NOR2_X2 U676 ( .A1(n606), .A2(n705), .ZN(n608) );
  INV_X1 U677 ( .A(KEYINPUT123), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(G54) );
  NAND2_X1 U679 ( .A1(n697), .A2(G472), .ZN(n610) );
  INV_X1 U680 ( .A(n705), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n613), .B(n612), .ZN(G36) );
  XNOR2_X1 U682 ( .A(n614), .B(G131), .ZN(G33) );
  NAND2_X1 U683 ( .A1(n697), .A2(G475), .ZN(n618) );
  XOR2_X1 U684 ( .A(KEYINPUT87), .B(KEYINPUT59), .Z(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U687 ( .A1(n619), .A2(n705), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n620), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U689 ( .A1(n697), .A2(G210), .ZN(n626) );
  XOR2_X1 U690 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT55), .B(KEYINPUT78), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U695 ( .A1(n627), .A2(n705), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U697 ( .A(G101), .B(n629), .Z(G3) );
  XOR2_X1 U698 ( .A(G104), .B(KEYINPUT111), .Z(n631) );
  NAND2_X1 U699 ( .A1(n632), .A2(n643), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n634) );
  NAND2_X1 U702 ( .A1(n632), .A2(n645), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(G107), .B(n635), .ZN(G9) );
  XNOR2_X1 U705 ( .A(G110), .B(n636), .ZN(G12) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U707 ( .A1(n345), .A2(n645), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(KEYINPUT112), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G45) );
  XOR2_X1 U711 ( .A(G146), .B(KEYINPUT113), .Z(n642) );
  NAND2_X1 U712 ( .A1(n345), .A2(n643), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n646), .A2(n643), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(G113), .ZN(G15) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U718 ( .A(G116), .B(n648), .ZN(G18) );
  XOR2_X1 U719 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n650) );
  XNOR2_X1 U720 ( .A(G125), .B(n347), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(G27) );
  XOR2_X1 U722 ( .A(G140), .B(n651), .Z(G42) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT117), .B(n656), .ZN(n661) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT118), .B(n659), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n662), .A2(n684), .ZN(n663) );
  XNOR2_X1 U730 ( .A(KEYINPUT119), .B(n663), .ZN(n680) );
  NAND2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U732 ( .A(n666), .B(KEYINPUT50), .Z(n671) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT49), .B(n669), .Z(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U738 ( .A(KEYINPUT51), .B(n676), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n686), .A2(n677), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT116), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n688) );
  INV_X1 U744 ( .A(n684), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n691), .B(KEYINPUT81), .ZN(n692) );
  NAND2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U750 ( .A1(G953), .A2(n694), .ZN(n696) );
  XNOR2_X1 U751 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n701), .A2(G478), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n705), .A2(n700), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n701), .A2(G217), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n705), .A2(n704), .ZN(G66) );
  XNOR2_X1 U759 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n720) );
  XNOR2_X1 U760 ( .A(G101), .B(n706), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n718) );
  NOR2_X1 U763 ( .A1(G953), .A2(n711), .ZN(n712) );
  XOR2_X1 U764 ( .A(KEYINPUT124), .B(n712), .Z(n716) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n722), .B(KEYINPUT127), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n721), .B(n727), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n731) );
  XNOR2_X1 U775 ( .A(n727), .B(G227), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G122), .B(n732), .ZN(G24) );
  XNOR2_X1 U780 ( .A(G137), .B(n733), .ZN(G39) );
  XNOR2_X1 U781 ( .A(G119), .B(n734), .ZN(G21) );
endmodule

