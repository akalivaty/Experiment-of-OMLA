

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n405), .B(n404), .Z(n565) );
  XNOR2_X1 U323 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U324 ( .A(n438), .B(n437), .ZN(n439) );
  NOR2_X1 U325 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U326 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U327 ( .A(n300), .B(n299), .ZN(n311) );
  XOR2_X1 U328 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n290) );
  XOR2_X1 U329 ( .A(G78GAT), .B(KEYINPUT22), .Z(n291) );
  INV_X1 U330 ( .A(KEYINPUT87), .ZN(n437) );
  NOR2_X1 U331 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U332 ( .A(n440), .B(n439), .ZN(n443) );
  XNOR2_X1 U333 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n487) );
  XNOR2_X1 U334 ( .A(n448), .B(KEYINPUT117), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n488), .B(n487), .ZN(n513) );
  XNOR2_X1 U336 ( .A(n461), .B(n290), .ZN(n564) );
  XOR2_X1 U337 ( .A(KEYINPUT36), .B(n537), .Z(n582) );
  XNOR2_X1 U338 ( .A(KEYINPUT79), .B(n409), .ZN(n537) );
  XOR2_X1 U339 ( .A(n466), .B(KEYINPUT28), .Z(n528) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  XOR2_X1 U343 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n293) );
  XNOR2_X1 U344 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U346 ( .A(n436), .B(n294), .Z(n300) );
  XOR2_X1 U347 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n295) );
  XOR2_X1 U349 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XOR2_X1 U351 ( .A(G92GAT), .B(G218GAT), .Z(n302) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n427) );
  XOR2_X1 U354 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n304) );
  XNOR2_X1 U355 ( .A(G99GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n370) );
  XOR2_X1 U357 ( .A(n427), .B(n370), .Z(n309) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n305), .B(KEYINPUT7), .ZN(n397) );
  XOR2_X1 U360 ( .A(G85GAT), .B(KEYINPUT77), .Z(n307) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n341) );
  XNOR2_X1 U363 ( .A(n397), .B(n341), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n550) );
  INV_X1 U366 ( .A(n550), .ZN(n409) );
  XOR2_X1 U367 ( .A(G99GAT), .B(G190GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U370 ( .A(G176GAT), .B(G71GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U373 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U374 ( .A(KEYINPUT84), .B(G120GAT), .Z(n319) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT85), .B(n320), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U379 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n324) );
  XNOR2_X1 U380 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U382 ( .A(n326), .B(n325), .Z(n331) );
  XNOR2_X1 U383 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n327), .B(KEYINPUT81), .ZN(n332) );
  XOR2_X1 U385 ( .A(G183GAT), .B(KEYINPUT18), .Z(n329) );
  XNOR2_X1 U386 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n418) );
  XNOR2_X1 U388 ( .A(n332), .B(n418), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n530) );
  XOR2_X1 U390 ( .A(G1GAT), .B(G127GAT), .Z(n351) );
  XOR2_X1 U391 ( .A(n332), .B(n351), .Z(n334) );
  NAND2_X1 U392 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n345) );
  XOR2_X1 U394 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n336) );
  XNOR2_X1 U395 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U397 ( .A(n337), .B(KEYINPUT4), .Z(n339) );
  XOR2_X1 U398 ( .A(G120GAT), .B(G57GAT), .Z(n368) );
  XNOR2_X1 U399 ( .A(G162GAT), .B(n368), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(n340), .B(KEYINPUT5), .Z(n343) );
  XNOR2_X1 U402 ( .A(n341), .B(KEYINPUT89), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U405 ( .A(KEYINPUT3), .B(G155GAT), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT2), .B(G148GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U408 ( .A(G141GAT), .B(n348), .ZN(n447) );
  XNOR2_X1 U409 ( .A(n349), .B(n447), .ZN(n465) );
  XNOR2_X1 U410 ( .A(KEYINPUT92), .B(n465), .ZN(n515) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G78GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n350), .B(KEYINPUT13), .ZN(n367) );
  XOR2_X1 U413 ( .A(n367), .B(n351), .Z(n353) );
  NAND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(n354), .B(KEYINPUT12), .Z(n357) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(G15GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n355), .B(KEYINPUT70), .ZN(n396) );
  XNOR2_X1 U419 ( .A(n396), .B(G64GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U421 ( .A(G57GAT), .B(G211GAT), .Z(n359) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(G155GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n361) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U427 ( .A(n363), .B(n362), .Z(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n484) );
  NOR2_X1 U429 ( .A1(n582), .A2(n484), .ZN(n366) );
  XNOR2_X1 U430 ( .A(KEYINPUT45), .B(n366), .ZN(n383) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(G176GAT), .B(G64GAT), .Z(n422) );
  XNOR2_X1 U433 ( .A(n369), .B(n422), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n370), .B(KEYINPUT32), .ZN(n372) );
  AND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U437 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U438 ( .A(G92GAT), .B(G85GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(G148GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U441 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n378) );
  XNOR2_X1 U442 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n569) );
  AND2_X1 U446 ( .A1(n383), .A2(n569), .ZN(n384) );
  XNOR2_X1 U447 ( .A(KEYINPUT113), .B(n384), .ZN(n406) );
  XOR2_X1 U448 ( .A(KEYINPUT29), .B(G1GAT), .Z(n386) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G113GAT), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n405) );
  XOR2_X1 U451 ( .A(G169GAT), .B(G8GAT), .Z(n417) );
  XOR2_X1 U452 ( .A(G141GAT), .B(G36GAT), .Z(n388) );
  XNOR2_X1 U453 ( .A(G50GAT), .B(G29GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n417), .B(n389), .Z(n391) );
  NAND2_X1 U456 ( .A1(G229GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n393) );
  XNOR2_X1 U459 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n398) );
  XOR2_X1 U462 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U463 ( .A1(n398), .A2(n399), .ZN(n403) );
  INV_X1 U464 ( .A(n398), .ZN(n401) );
  INV_X1 U465 ( .A(n399), .ZN(n400) );
  NAND2_X1 U466 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U468 ( .A1(n406), .A2(n565), .ZN(n415) );
  XNOR2_X1 U469 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n569), .B(KEYINPUT41), .ZN(n557) );
  NAND2_X1 U471 ( .A1(n565), .A2(n557), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n407), .B(KEYINPUT46), .ZN(n408) );
  AND2_X1 U473 ( .A1(n484), .A2(n408), .ZN(n410) );
  AND2_X1 U474 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n413), .B(KEYINPUT47), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT48), .ZN(n525) );
  XOR2_X1 U479 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n421), .B(KEYINPUT93), .Z(n424) );
  XNOR2_X1 U483 ( .A(n422), .B(KEYINPUT94), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U485 ( .A(G204GAT), .B(G211GAT), .Z(n426) );
  XNOR2_X1 U486 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n441) );
  XOR2_X1 U488 ( .A(n441), .B(n427), .Z(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n460) );
  NOR2_X1 U490 ( .A1(n525), .A2(n460), .ZN(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT54), .B(n430), .Z(n431) );
  NOR2_X1 U492 ( .A1(n515), .A2(n431), .ZN(n563) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U494 ( .A(G22GAT), .B(KEYINPUT88), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n445) );
  XNOR2_X1 U496 ( .A(G218GAT), .B(G106GAT), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n291), .B(n434), .ZN(n435) );
  XOR2_X1 U498 ( .A(n436), .B(n435), .Z(n440) );
  NAND2_X1 U499 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n441), .B(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n466) );
  AND2_X1 U504 ( .A1(n563), .A2(n466), .ZN(n450) );
  INV_X1 U505 ( .A(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U506 ( .A1(n530), .A2(n451), .ZN(n560) );
  NAND2_X1 U507 ( .A1(n537), .A2(n560), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n475) );
  NAND2_X1 U509 ( .A1(n569), .A2(n565), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT75), .ZN(n489) );
  NOR2_X1 U511 ( .A1(n537), .A2(n484), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT16), .B(n455), .ZN(n472) );
  INV_X1 U513 ( .A(n530), .ZN(n519) );
  INV_X1 U514 ( .A(n460), .ZN(n517) );
  NAND2_X1 U515 ( .A1(n519), .A2(n517), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n456), .A2(n466), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT96), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT27), .B(n460), .Z(n467) );
  NOR2_X1 U521 ( .A1(n466), .A2(n519), .ZN(n461) );
  AND2_X1 U522 ( .A1(n467), .A2(n564), .ZN(n462) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n470) );
  OR2_X1 U524 ( .A1(n519), .A2(n528), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n515), .A2(n467), .ZN(n526) );
  NOR2_X1 U526 ( .A1(n468), .A2(n526), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n471), .Z(n486) );
  AND2_X1 U528 ( .A1(n472), .A2(n486), .ZN(n504) );
  NAND2_X1 U529 ( .A1(n489), .A2(n504), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(n473), .ZN(n481) );
  NAND2_X1 U531 ( .A1(n481), .A2(n515), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n476), .Z(G1324GAT) );
  XOR2_X1 U534 ( .A(G8GAT), .B(KEYINPUT101), .Z(n478) );
  NAND2_X1 U535 ( .A1(n481), .A2(n517), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U538 ( .A1(n481), .A2(n519), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n481), .A2(n528), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  INV_X1 U543 ( .A(n484), .ZN(n574) );
  NOR2_X1 U544 ( .A1(n582), .A2(n574), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n513), .A2(n489), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT105), .B(n491), .ZN(n500) );
  NAND2_X1 U549 ( .A1(n500), .A2(n515), .ZN(n494) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n500), .A2(n517), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT107), .ZN(n499) );
  NAND2_X1 U556 ( .A1(n500), .A2(n519), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1330GAT) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n502) );
  NAND2_X1 U561 ( .A1(n528), .A2(n500), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n557), .ZN(n503) );
  NOR2_X1 U564 ( .A1(n565), .A2(n503), .ZN(n512) );
  AND2_X1 U565 ( .A1(n512), .A2(n504), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n515), .A2(n509), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n505), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n517), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n519), .A2(n509), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U574 ( .A1(n509), .A2(n528), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT109), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n521), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n523) );
  NAND2_X1 U585 ( .A1(n521), .A2(n528), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U589 ( .A(n527), .B(KEYINPUT114), .Z(n541) );
  OR2_X1 U590 ( .A1(n541), .A2(n528), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n538), .A2(n565), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U595 ( .A1(n538), .A2(n557), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  NAND2_X1 U598 ( .A1(n538), .A2(n574), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  INV_X1 U604 ( .A(n564), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n565), .A2(n549), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U609 ( .A1(n549), .A2(n557), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n549), .A2(n574), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT116), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n565), .A2(n560), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n574), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n581) );
  INV_X1 U631 ( .A(n581), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n581), .A2(n569), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

