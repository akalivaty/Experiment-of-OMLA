//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n205), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(new_n205), .C1(new_n210), .C2(new_n216), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n213), .A2(new_n227), .A3(new_n215), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n210), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(KEYINPUT25), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n218), .A2(new_n220), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n236));
  INV_X1    g035(.A(G134gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G127gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(G127gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT69), .B(G134gat), .Z(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n242), .B2(G127gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT68), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(KEYINPUT26), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n206), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n222), .A2(G183gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT27), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT28), .B1(new_n258), .B2(new_n221), .ZN(new_n259));
  AND2_X1   g058(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT28), .B(new_n221), .C1(new_n260), .C2(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT28), .A4(new_n221), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n212), .B(new_n252), .C1(new_n259), .C2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n233), .A2(new_n246), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n246), .B1(new_n233), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n204), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT71), .B(new_n204), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n233), .A2(new_n267), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n245), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n233), .A2(new_n246), .A3(new_n267), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT71), .B1(new_n284), .B2(new_n204), .ZN(new_n285));
  INV_X1    g084(.A(new_n273), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT32), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(new_n203), .A3(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT34), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT34), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n282), .A2(new_n290), .A3(new_n203), .A4(new_n283), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n291), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(KEYINPUT32), .B2(new_n274), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n280), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n292), .ZN(new_n297));
  INV_X1    g096(.A(new_n279), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n274), .B2(new_n275), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(new_n294), .A3(KEYINPUT32), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT85), .Z(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT77), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306));
  AND2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  OAI22_X1  g107(.A1(new_n305), .A2(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT76), .B1(new_n311), .B2(G141gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(G141gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n311), .A2(G141gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n307), .A2(new_n308), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n310), .A2(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT22), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  INV_X1    g129(.A(G218gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n328), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n329), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n323), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G204gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G197gat), .ZN(new_n341));
  INV_X1    g140(.A(G197gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G204gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n328), .B(new_n332), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G141gat), .B(G148gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n321), .B1(new_n349), .B2(KEYINPUT2), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n350), .B(new_n338), .C1(new_n351), .C2(new_n309), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n352), .B2(new_n323), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n303), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR3_X1    g155(.A1(new_n339), .A2(new_n353), .A3(new_n302), .ZN(new_n357));
  OAI211_X1 g156(.A(KEYINPUT86), .B(new_n303), .C1(new_n339), .C2(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G78gat), .B(G106gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT84), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G22gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n362), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n364), .B2(new_n367), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT87), .B(G50gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n364), .A2(new_n367), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n365), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n371), .B1(new_n375), .B2(new_n368), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n296), .B(new_n301), .C1(new_n373), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT73), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n233), .A2(new_n379), .A3(new_n267), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n233), .A2(new_n267), .B1(new_n323), .B2(new_n379), .ZN(new_n382));
  INV_X1    g181(.A(new_n348), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n323), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n281), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n348), .B1(new_n386), .B2(new_n380), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  INV_X1    g188(.A(G64gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n384), .B2(new_n387), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n383), .B1(new_n381), .B2(new_n382), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n386), .A2(new_n348), .A3(new_n380), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n394), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n395), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n350), .B1(new_n351), .B2(new_n309), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n245), .A3(new_n352), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT78), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(new_n245), .A3(new_n410), .A4(new_n352), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT4), .B1(new_n245), .B2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT69), .B(G134gat), .ZN(new_n416));
  INV_X1    g215(.A(G127gat), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n239), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(KEYINPUT1), .B2(new_n234), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n322), .A2(new_n419), .A3(new_n420), .A4(new_n241), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n421), .A2(new_n415), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n412), .A2(new_n413), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n245), .B(new_n406), .ZN(new_n426));
  INV_X1    g225(.A(new_n413), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n409), .A2(new_n411), .B1(new_n421), .B2(new_n414), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n425), .A3(new_n413), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G1gat), .B(G29gat), .Z(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n405), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n437), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n439), .A3(new_n431), .ZN(new_n440));
  INV_X1    g239(.A(new_n404), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n439), .B1(new_n429), .B2(new_n431), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n441), .B(new_n440), .C1(new_n444), .C2(new_n405), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT30), .A4(new_n394), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT75), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n403), .A2(new_n443), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n202), .B1(new_n377), .B2(new_n449), .ZN(new_n450));
  AND4_X1   g249(.A1(new_n445), .A2(new_n403), .A3(new_n443), .A4(new_n448), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n299), .B1(new_n297), .B2(new_n300), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n372), .B1(new_n369), .B2(new_n370), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n375), .A2(new_n371), .A3(new_n368), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n451), .A2(KEYINPUT35), .A3(new_n454), .A4(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n452), .B2(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n296), .A2(KEYINPUT36), .A3(new_n301), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n373), .A2(new_n376), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n449), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n445), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n394), .B1(new_n388), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n468), .C1(new_n466), .C2(new_n388), .ZN(new_n469));
  INV_X1    g268(.A(new_n388), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n393), .B1(new_n470), .B2(KEYINPUT37), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n397), .B2(new_n400), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT38), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n465), .A2(new_n395), .A3(new_n469), .A4(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n426), .A2(new_n427), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(KEYINPUT39), .C1(new_n430), .C2(new_n413), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n414), .A2(new_n421), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n412), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n427), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n480), .A3(new_n439), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n481), .A2(KEYINPUT88), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n481), .B2(KEYINPUT88), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n483), .A2(new_n484), .A3(new_n444), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n403), .A2(new_n448), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n474), .A2(new_n487), .A3(new_n457), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n464), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n459), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n390), .B2(G57gat), .ZN(new_n492));
  INV_X1    g291(.A(G57gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n492), .B(new_n494), .C1(new_n493), .C2(G64gat), .ZN(new_n495));
  INV_X1    g294(.A(G71gat), .ZN(new_n496));
  INV_X1    g295(.A(G78gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT9), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n493), .A2(G64gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n390), .A2(G57gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT9), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G71gat), .B(G78gat), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n499), .A2(new_n495), .B1(new_n503), .B2(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT96), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G127gat), .B(G155gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n330), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G8gat), .ZN(new_n523));
  OAI21_X1  g322(.A(G183gat), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n224), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G231gat), .ZN(new_n528));
  INV_X1    g327(.A(G233gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n524), .B2(new_n527), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n517), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n532), .A2(new_n533), .A3(new_n517), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n515), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n514), .A3(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n392), .ZN(new_n543));
  NAND2_X1  g342(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n542), .B2(new_n392), .ZN(new_n545));
  NAND4_X1  g344(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G99gat), .ZN(new_n548));
  INV_X1    g347(.A(G106gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n541), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n543), .A2(new_n552), .A3(new_n545), .A4(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G43gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(G50gat), .ZN(new_n559));
  INV_X1    g358(.A(G50gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(G43gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT91), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT15), .ZN(new_n563));
  INV_X1    g362(.A(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT14), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(new_n568), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n572), .B2(new_n569), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT92), .B1(new_n573), .B2(KEYINPUT17), .ZN(new_n574));
  INV_X1    g373(.A(new_n570), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n569), .B1(new_n563), .B2(new_n571), .ZN(new_n576));
  OAI211_X1 g375(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI221_X1 g377(.A(new_n554), .B1(KEYINPUT17), .B2(new_n573), .C1(new_n574), .C2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT41), .ZN(new_n581));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT97), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n573), .A2(new_n554), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n580), .B1(new_n579), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT99), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n580), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n554), .B1(new_n574), .B2(new_n578), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n573), .A2(KEYINPUT17), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n592), .B2(new_n584), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n583), .A2(new_n581), .ZN(new_n597));
  XOR2_X1   g396(.A(G134gat), .B(G162gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n588), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n540), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT100), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n540), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n490), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n575), .A2(new_n576), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n523), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n574), .B2(new_n578), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT93), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n523), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT18), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n526), .A2(new_n573), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(KEYINPUT94), .A3(new_n615), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n614), .B(KEYINPUT13), .Z(new_n621));
  OR3_X1    g420(.A1(new_n609), .A2(new_n523), .A3(KEYINPUT94), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n612), .A2(KEYINPUT18), .A3(new_n614), .A4(new_n615), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT90), .ZN(new_n627));
  XOR2_X1   g426(.A(G113gat), .B(G141gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G169gat), .B(G197gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n632), .A2(new_n618), .A3(new_n623), .A4(new_n624), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT101), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n500), .A2(KEYINPUT96), .A3(new_n505), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT96), .B1(new_n500), .B2(new_n505), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n554), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n551), .A2(new_n553), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n506), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT10), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(KEYINPUT10), .C1(new_n640), .C2(new_n641), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n639), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n554), .A2(new_n509), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n511), .B2(new_n554), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n638), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n248), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n340), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n608), .A2(new_n636), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n465), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(G8gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n486), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n486), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(G8gat), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n665), .B1(new_n668), .B2(new_n664), .ZN(G1325gat));
  AOI21_X1  g468(.A(G15gat), .B1(new_n659), .B2(new_n454), .ZN(new_n670));
  INV_X1    g469(.A(new_n461), .ZN(new_n671));
  INV_X1    g470(.A(new_n462), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n659), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n463), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n603), .A2(KEYINPUT105), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n601), .A2(new_n680), .A3(new_n602), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI211_X1 g481(.A(KEYINPUT44), .B(new_n682), .C1(new_n459), .C2(new_n489), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n603), .B1(new_n459), .B2(new_n489), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(KEYINPUT104), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  INV_X1    g487(.A(new_n603), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n464), .A2(new_n488), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n450), .A2(new_n458), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n692), .B2(KEYINPUT44), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n684), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n540), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n636), .A2(new_n658), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n465), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n692), .A2(new_n697), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n564), .A3(new_n465), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(new_n486), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n699), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n565), .A3(new_n486), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n685), .B2(new_n686), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n692), .A2(new_n688), .A3(KEYINPUT44), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n683), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n697), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n565), .B1(new_n717), .B2(new_n486), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n712), .A2(new_n711), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n717), .A2(G43gat), .A3(new_n673), .ZN(new_n722));
  AOI21_X1  g521(.A(G43gat), .B1(new_n702), .B2(new_n454), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT47), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n727), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n699), .B2(new_n457), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n702), .A2(new_n560), .A3(new_n463), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(KEYINPUT48), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n560), .B1(new_n717), .B2(new_n463), .ZN(new_n735));
  INV_X1    g534(.A(new_n731), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n634), .A2(new_n635), .ZN(new_n739));
  INV_X1    g538(.A(new_n658), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n608), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n465), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  INV_X1    g542(.A(new_n741), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n486), .B(new_n745), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n744), .A2(new_n746), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n746), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT49), .B(G64gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n741), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT109), .B(KEYINPUT110), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1333gat));
  INV_X1    g552(.A(new_n454), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n496), .B1(new_n744), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n741), .A2(G71gat), .A3(new_n673), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n463), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n540), .A2(new_n739), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n694), .A2(new_n658), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT111), .B1(new_n762), .B2(new_n700), .ZN(new_n763));
  INV_X1    g562(.A(new_n761), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n716), .A2(new_n740), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n465), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n767), .A3(G85gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(new_n692), .B2(KEYINPUT112), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n685), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n769), .B2(new_n771), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT113), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT113), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n465), .A2(new_n542), .A3(new_n658), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT114), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n768), .A2(new_n779), .ZN(G1336gat));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(G92gat), .C1(new_n762), .C2(new_n746), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n761), .B1(new_n685), .B2(new_n770), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n692), .A2(KEYINPUT112), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n740), .B1(new_n786), .B2(new_n772), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n746), .A2(G92gat), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n787), .A2(new_n788), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n788), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n740), .B(new_n791), .C1(new_n786), .C2(new_n772), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n694), .A2(new_n658), .A3(new_n486), .A4(new_n761), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(KEYINPUT115), .B1(new_n793), .B2(G92gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n794), .B2(new_n781), .ZN(G1337gat));
  INV_X1    g594(.A(new_n673), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n762), .A2(new_n548), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n754), .A2(new_n740), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n775), .A2(new_n776), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n548), .ZN(G1338gat));
  NOR2_X1   g599(.A1(new_n457), .A2(G106gat), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n658), .B(new_n801), .C1(new_n773), .C2(new_n774), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n716), .A2(new_n740), .A3(new_n457), .A4(new_n764), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n549), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT53), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n802), .B(new_n806), .C1(new_n803), .C2(new_n549), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1339gat));
  AOI21_X1  g607(.A(new_n614), .B1(new_n612), .B2(new_n615), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n631), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n635), .A2(new_n658), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n638), .B(new_n646), .C1(new_n650), .C2(KEYINPUT10), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n648), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n815), .B(new_n639), .C1(new_n645), .C2(new_n647), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n655), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n656), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n648), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n655), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT116), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n812), .B1(new_n636), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT117), .B(new_n812), .C1(new_n636), .C2(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n682), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n635), .A2(new_n811), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n679), .A2(new_n681), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n540), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n739), .A2(new_n658), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n605), .A2(new_n607), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n377), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n465), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n748), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n636), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n636), .A2(G113gat), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT118), .Z(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n843), .B2(new_n846), .ZN(G1340gat));
  NAND2_X1  g646(.A1(new_n842), .A2(new_n658), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n540), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(G127gat), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n843), .B2(new_n603), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n689), .A2(new_n707), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT119), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n841), .A2(new_n416), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n673), .A2(new_n700), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n746), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n739), .A2(new_n818), .A3(new_n822), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n812), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n603), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n540), .B1(new_n864), .B2(new_n834), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n463), .B1(new_n838), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n463), .B1(new_n835), .B2(new_n838), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(KEYINPUT57), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n636), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n463), .B(new_n860), .C1(new_n835), .C2(new_n838), .ZN(new_n871));
  OR4_X1    g670(.A1(G141gat), .A2(new_n871), .A3(new_n636), .A4(new_n748), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT120), .B(KEYINPUT58), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n874));
  NAND2_X1  g673(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n874), .A2(new_n870), .A3(new_n872), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n873), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(G148gat), .C1(new_n869), .C2(new_n740), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n861), .A2(new_n740), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n837), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n689), .B1(new_n812), .B2(new_n862), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n603), .A2(new_n832), .A3(new_n826), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n695), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n605), .A2(KEYINPUT121), .A3(new_n607), .A4(new_n836), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n463), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n880), .A2(new_n881), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G148gat), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT122), .B1(new_n892), .B2(KEYINPUT59), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n894), .B(new_n878), .C1(new_n891), .C2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n879), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OR4_X1    g695(.A1(G148gat), .A2(new_n868), .A3(new_n740), .A4(new_n861), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1345gat));
  INV_X1    g697(.A(new_n869), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(G155gat), .A3(new_n540), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n871), .A2(new_n695), .A3(new_n748), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(G155gat), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(G1346gat));
  XOR2_X1   g702(.A(KEYINPUT77), .B(G162gat), .Z(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n869), .B2(new_n682), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n854), .A2(new_n904), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n871), .B2(new_n906), .ZN(G1347gat));
  OAI21_X1  g706(.A(KEYINPUT123), .B1(new_n839), .B2(new_n465), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(new_n700), .C1(new_n835), .C2(new_n838), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n377), .B(new_n746), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n247), .A3(new_n739), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n707), .A2(new_n465), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n840), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n636), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(G1348gat));
  NOR3_X1   g715(.A1(new_n914), .A2(new_n248), .A3(new_n740), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n658), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n248), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n908), .A2(new_n910), .ZN(new_n920));
  INV_X1    g719(.A(new_n377), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n540), .A2(new_n263), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n748), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n223), .A2(new_n225), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n914), .B2(new_n695), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT124), .B(KEYINPUT60), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  OR2_X1    g725(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n927));
  NAND2_X1  g726(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n927), .A2(new_n923), .A3(new_n928), .A4(new_n925), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n926), .A2(new_n929), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n914), .B2(new_n603), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  INV_X1    g731(.A(new_n682), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n221), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1351gat));
  NAND4_X1  g734(.A1(new_n880), .A2(new_n796), .A3(new_n890), .A4(new_n913), .ZN(new_n936));
  OAI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n636), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n457), .B1(new_n908), .B2(new_n910), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(new_n748), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n342), .A3(new_n796), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n940), .B2(new_n636), .ZN(G1352gat));
  XNOR2_X1  g740(.A(KEYINPUT125), .B(G204gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n740), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n938), .A2(new_n796), .A3(new_n748), .A4(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n936), .A2(KEYINPUT126), .A3(new_n740), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT126), .B1(new_n936), .B2(new_n740), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(G1353gat));
  NAND4_X1  g749(.A1(new_n939), .A2(new_n330), .A3(new_n540), .A4(new_n796), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n936), .A2(new_n695), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT63), .B(G211gat), .C1(new_n936), .C2(new_n695), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n953), .B2(new_n955), .ZN(G1354gat));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n331), .A3(new_n796), .A4(new_n933), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n936), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n936), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n603), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n331), .ZN(G1355gat));
endmodule


