//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(KEYINPUT87), .A2(G143), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND4_X1  g003(.A1(new_n187), .A2(G214), .A3(new_n188), .A4(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT87), .B(G143), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT18), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(G125), .A2(G140), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n190), .B(G131), .C1(new_n191), .C2(new_n192), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n196), .B(new_n206), .C1(new_n194), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n193), .A2(new_n195), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n207), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n207), .A2(new_n210), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(KEYINPUT91), .A3(new_n210), .A4(new_n207), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  OAI211_X1 g033(.A(G146), .B(new_n218), .C1(new_n201), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n199), .B2(new_n200), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n204), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n208), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT89), .B(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(G475), .A2(G902), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT19), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n203), .B(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n220), .B1(new_n234), .B2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT88), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n220), .C1(new_n234), .C2(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n209), .A2(new_n207), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n208), .A3(new_n229), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n232), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT20), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n231), .A2(new_n244), .A3(new_n232), .A4(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n229), .A2(KEYINPUT92), .ZN(new_n247));
  AOI21_X1  g061(.A(G902), .B1(new_n226), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n226), .B2(new_n247), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G475), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT73), .B(G902), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT94), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT94), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G122), .ZN(new_n266));
  INV_X1    g080(.A(G122), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G116), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G107), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n254), .A2(G143), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n255), .B1(new_n272), .B2(KEYINPUT13), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n264), .B(new_n271), .C1(new_n278), .C2(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n270), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT95), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT14), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n268), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT96), .B1(new_n283), .B2(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n268), .A2(new_n282), .ZN(new_n285));
  INV_X1    g099(.A(new_n266), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n286), .B(new_n287), .C1(new_n282), .C2(new_n268), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G107), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n260), .A2(G134), .A3(new_n261), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n264), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n281), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(G217), .A3(new_n189), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n279), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n279), .B2(new_n293), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n253), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n301));
  OAI21_X1  g115(.A(G478), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n303), .A2(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n301), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G952), .ZN(new_n310));
  AOI211_X1 g124(.A(G953), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n311));
  AOI211_X1 g125(.A(new_n189), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT21), .B(G898), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n251), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G221), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n294), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n189), .A2(G227), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n322), .B(new_n323), .Z(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n325), .B(new_n326), .C1(new_n327), .C2(G107), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n270), .B(G104), .C1(KEYINPUT77), .C2(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n325), .A2(new_n326), .B1(new_n270), .B2(G104), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n330), .B2(new_n332), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n331), .B1(new_n328), .B2(new_n329), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n336), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n204), .A2(G143), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n256), .A2(G146), .ZN(new_n344));
  OAI21_X1  g158(.A(G128), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n256), .A2(G146), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n204), .A2(G143), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n254), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(KEYINPUT0), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT0), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n337), .A2(new_n338), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n330), .A2(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n339), .A2(new_n333), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G101), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n340), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n342), .A2(new_n354), .A3(new_n355), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT1), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT65), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G143), .B(G146), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n254), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n346), .A2(new_n347), .A3(new_n254), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n369), .A2(new_n370), .B1(new_n346), .B2(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n327), .A2(G107), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n270), .A2(G104), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n336), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n339), .B2(new_n336), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n375), .A3(KEYINPUT10), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n380));
  OAI21_X1  g194(.A(G128), .B1(new_n350), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n381), .A2(new_n348), .B1(KEYINPUT1), .B2(new_n343), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(KEYINPUT10), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n362), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G137), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT64), .B1(new_n386), .B2(G134), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n263), .A3(G137), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT11), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n263), .B2(G137), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(KEYINPUT11), .A3(G134), .ZN(new_n393));
  AND4_X1   g207(.A1(new_n195), .A2(new_n390), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n195), .B1(new_n395), .B2(new_n390), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n362), .A2(new_n378), .A3(new_n397), .A4(new_n384), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n324), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n371), .A2(new_n375), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n398), .B1(new_n383), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT12), .B(new_n398), .C1(new_n383), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n400), .A2(new_n407), .A3(new_n324), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n321), .B(new_n253), .C1(new_n401), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(G469), .A2(G902), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n399), .A2(new_n400), .A3(new_n324), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n407), .ZN(new_n412));
  INV_X1    g226(.A(new_n324), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n409), .B(new_n410), .C1(new_n321), .C2(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n316), .A2(new_n320), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n352), .B(new_n349), .C1(new_n394), .C2(new_n396), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n395), .A2(new_n195), .A3(new_n390), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n263), .A2(G137), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n386), .A2(G134), .ZN(new_n422));
  OAI21_X1  g236(.A(G131), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n367), .A2(new_n368), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n370), .B1(new_n424), .B2(G128), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n367), .A2(new_n346), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n420), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G116), .B(G119), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT2), .B(G113), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n419), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT28), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT28), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n418), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT72), .B1(new_n431), .B2(new_n435), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(G101), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(KEYINPUT29), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n396), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n353), .B1(new_n449), .B2(new_n420), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n420), .A2(new_n423), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n426), .B1(new_n381), .B2(new_n348), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT30), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n419), .A2(new_n427), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n430), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n446), .B(new_n445), .C1(new_n457), .C2(new_n432), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n445), .A2(KEYINPUT70), .A3(new_n446), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT70), .B1(new_n445), .B2(new_n446), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n434), .A2(new_n436), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n458), .A2(new_n462), .A3(new_n466), .A4(new_n463), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n448), .A2(new_n465), .A3(new_n253), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G472), .ZN(new_n469));
  NOR2_X1   g283(.A1(G472), .A2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n431), .A2(new_n473), .A3(new_n447), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n431), .B2(new_n447), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n457), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT31), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n430), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n419), .A2(new_n427), .A3(new_n455), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n455), .B1(new_n419), .B2(new_n427), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n431), .A2(new_n447), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT67), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n431), .A2(new_n473), .A3(new_n447), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n461), .B1(new_n434), .B2(new_n436), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n482), .A2(new_n484), .A3(new_n477), .A4(new_n485), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT69), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n474), .A2(new_n475), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n477), .A4(new_n482), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n471), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT32), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(KEYINPUT32), .B(new_n471), .C1(new_n488), .C2(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n469), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G119), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G128), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n254), .A2(G119), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n501), .A2(G128), .ZN(new_n509));
  AND2_X1   g323(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n511), .A3(KEYINPUT75), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(G110), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n508), .A2(new_n509), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT24), .B(G110), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n223), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G110), .B1(new_n507), .B2(new_n511), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n220), .B(new_n205), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT22), .B(G137), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n523), .A3(new_n527), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n253), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT25), .ZN(new_n532));
  INV_X1    g346(.A(G217), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n253), .B2(G234), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n529), .A2(new_n535), .A3(new_n253), .A4(new_n530), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n532), .A2(new_n539), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n529), .A2(new_n530), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n534), .A2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G214), .B1(G237), .B2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G210), .B1(G237), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n353), .A2(G125), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n353), .A2(KEYINPUT83), .A3(G125), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(KEYINPUT84), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT84), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT83), .B1(new_n353), .B2(G125), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n551), .B(new_n197), .C1(new_n349), .C2(new_n352), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n452), .A2(new_n197), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G224), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT85), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n560), .B(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n342), .A2(new_n355), .A3(new_n361), .A4(new_n479), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n265), .A2(G119), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G113), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n428), .B2(new_n566), .ZN(new_n570));
  INV_X1    g384(.A(new_n429), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n428), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n375), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G122), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n565), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(KEYINPUT82), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n565), .B2(new_n573), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT6), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n578), .A2(KEYINPUT6), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n564), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n565), .A2(new_n573), .A3(new_n574), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n379), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n574), .B(KEYINPUT8), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n569), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n428), .B2(new_n571), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n583), .B(new_n584), .C1(new_n379), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n552), .A2(new_n559), .A3(new_n553), .ZN(new_n590));
  OR2_X1    g404(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g405(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n563), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n554), .A2(new_n558), .A3(new_n563), .A4(new_n559), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT7), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n318), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n549), .B1(new_n581), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n582), .A2(new_n588), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n578), .A2(KEYINPUT6), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n565), .A2(new_n573), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n582), .B1(new_n604), .B2(new_n577), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n605), .B2(KEYINPUT6), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n548), .B(new_n602), .C1(new_n606), .C2(new_n564), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n547), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n417), .A2(new_n500), .A3(new_n545), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n299), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n613));
  OR3_X1    g427(.A1(new_n297), .A2(new_n298), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  OAI22_X1  g429(.A1(new_n297), .A2(new_n298), .B1(KEYINPUT99), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n614), .A2(G478), .A3(new_n253), .A4(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n246), .A2(new_n250), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT100), .Z(new_n619));
  INV_X1    g433(.A(new_n315), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n608), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n416), .A2(new_n320), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n252), .B1(new_n488), .B2(new_n495), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n496), .B1(new_n624), .B2(G472), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n625), .A3(new_n545), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n245), .A2(KEYINPUT101), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n243), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n242), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n634), .A2(new_n250), .ZN(new_n635));
  AND4_X1   g449(.A1(new_n309), .A2(new_n608), .A3(new_n620), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n524), .B(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n643), .B2(new_n543), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n524), .B1(KEYINPUT36), .B2(new_n528), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n520), .A2(new_n523), .A3(new_n642), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n641), .A2(new_n645), .A3(new_n543), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n538), .A2(new_n540), .A3(new_n648), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n547), .B(new_n649), .C1(new_n599), .C2(new_n607), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n417), .A2(new_n625), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G110), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  NAND3_X1  g468(.A1(new_n500), .A2(new_n650), .A3(new_n622), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n311), .B1(new_n312), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n634), .A2(new_n309), .A3(new_n250), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT106), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n416), .A2(new_n320), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n491), .A2(new_n494), .ZN(new_n664));
  INV_X1    g478(.A(new_n489), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n486), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT68), .B1(new_n486), .B2(KEYINPUT31), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n470), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT32), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n496), .A2(new_n497), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n663), .B1(new_n673), .B2(new_n469), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n659), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .A4(new_n650), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n662), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XNOR2_X1  g493(.A(new_n657), .B(KEYINPUT39), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n622), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT108), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n599), .A2(new_n607), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n251), .A2(new_n309), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n432), .A2(new_n433), .ZN(new_n690));
  INV_X1    g504(.A(new_n461), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n476), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n692), .B2(G902), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n689), .B1(new_n673), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n688), .A2(new_n546), .A3(new_n649), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n256), .ZN(G45));
  AND2_X1   g511(.A1(new_n618), .A2(new_n658), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n500), .A2(new_n650), .A3(new_n622), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  OAI21_X1  g514(.A(new_n253), .B1(new_n401), .B2(new_n408), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n409), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n701), .A2(KEYINPUT109), .A3(G469), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n319), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n500), .A2(new_n706), .A3(new_n545), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n621), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT41), .B(G113), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  INV_X1    g524(.A(new_n545), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n673), .B2(new_n469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n636), .A3(new_n706), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  INV_X1    g528(.A(new_n649), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n316), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n500), .A2(new_n716), .A3(new_n706), .A4(new_n608), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT110), .B(G119), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G21));
  AOI211_X1 g533(.A(new_n547), .B(new_n689), .C1(new_n599), .C2(new_n607), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n486), .A2(KEYINPUT31), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n691), .B1(new_n437), .B2(new_n438), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n664), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n470), .ZN(new_n724));
  INV_X1    g538(.A(G472), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n724), .B1(new_n623), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n315), .A3(new_n711), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n720), .A2(new_n727), .A3(new_n706), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  OAI211_X1 g543(.A(new_n724), .B(new_n618), .C1(new_n623), .C2(new_n725), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n649), .A2(new_n657), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n706), .A2(new_n731), .A3(new_n608), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n498), .B2(new_n499), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n671), .A2(KEYINPUT111), .A3(new_n672), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n469), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n663), .A2(new_n547), .A3(new_n685), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n545), .A4(new_n698), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n712), .A2(new_n742), .A3(new_n739), .A4(new_n698), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n195), .ZN(G33));
  NAND3_X1  g559(.A1(new_n712), .A2(new_n675), .A3(new_n739), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NOR2_X1   g561(.A1(new_n685), .A2(new_n547), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n409), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n415), .B(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n410), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n320), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n680), .ZN(new_n758));
  INV_X1    g572(.A(new_n625), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n617), .A2(new_n612), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n246), .A3(new_n250), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n761), .B1(KEYINPUT112), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(new_n715), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n758), .B1(KEYINPUT44), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n749), .B(new_n768), .C1(KEYINPUT44), .C2(new_n767), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n386), .ZN(G39));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n757), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n757), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n749), .A2(new_n500), .A3(new_n545), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n698), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT114), .B(G140), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G42));
  NAND3_X1  g594(.A1(new_n673), .A2(new_n311), .A3(new_n693), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n545), .A3(new_n706), .A4(new_n748), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT121), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT121), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n619), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(G952), .A3(new_n189), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT48), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n765), .A2(new_n311), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n706), .A3(new_n748), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n738), .A2(new_n545), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n788), .A2(KEYINPUT48), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n787), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n251), .A2(new_n760), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n784), .A2(new_n785), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n726), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n791), .A2(new_n715), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n706), .A2(new_n547), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n688), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n790), .A2(new_n799), .A3(new_n545), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n802), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n704), .A2(new_n705), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n319), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n773), .B2(new_n775), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n748), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n808), .A2(new_n802), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n812), .B1(new_n818), .B2(new_n809), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n796), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n811), .B(new_n801), .C1(new_n823), .C2(new_n810), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n824), .B2(KEYINPUT51), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n819), .A2(KEYINPUT122), .A3(new_n820), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n810), .A2(new_n608), .A3(new_n706), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n699), .A2(new_n733), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n673), .A2(new_n693), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n657), .B(KEYINPUT117), .Z(new_n832));
  NOR2_X1   g646(.A1(new_n663), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n720), .A3(new_n649), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n678), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n662), .B2(new_n677), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n713), .A2(new_n717), .A3(new_n728), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n609), .B(new_n651), .C1(new_n621), .C2(new_n707), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n251), .A2(new_n308), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n608), .A2(new_n620), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n608), .A2(new_n620), .A3(new_n618), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n608), .A2(KEYINPUT116), .A3(new_n620), .A4(new_n844), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n608), .A2(KEYINPUT115), .A3(new_n620), .A4(new_n618), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n630), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n500), .A2(new_n308), .A3(new_n635), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n732), .B(new_n739), .C1(new_n856), .C2(new_n731), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n741), .A2(new_n857), .A3(new_n743), .A4(new_n746), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n847), .A2(new_n851), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n850), .A2(new_n852), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n626), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n713), .A2(new_n717), .A3(new_n728), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n842), .A3(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n741), .A2(new_n857), .A3(new_n743), .A4(new_n746), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND4_X1   g681(.A1(KEYINPUT52), .A2(new_n678), .A3(new_n830), .A4(new_n834), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n838), .B2(new_n834), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT118), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n837), .A2(new_n871), .A3(new_n839), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n860), .B1(new_n873), .B2(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n868), .A2(new_n869), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n867), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT118), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n871), .B1(new_n837), .B2(new_n839), .ZN(new_n882));
  OAI211_X1 g696(.A(KEYINPUT53), .B(new_n859), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .A3(new_n876), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n880), .A2(new_n883), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n827), .A2(new_n828), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(G952), .B2(G953), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n813), .B(KEYINPUT49), .Z(new_n891));
  NOR4_X1   g705(.A1(new_n891), .A2(new_n547), .A3(new_n831), .A4(new_n761), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n320), .A3(new_n545), .A4(new_n687), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(G75));
  AOI211_X1 g708(.A(new_n879), .B(KEYINPUT53), .C1(new_n840), .C2(new_n859), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT119), .B1(new_n885), .B2(new_n876), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n253), .B1(new_n897), .B2(new_n883), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n549), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n606), .B(new_n564), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n903), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n189), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n410), .B(KEYINPUT57), .Z(new_n908));
  AOI21_X1  g722(.A(new_n884), .B1(new_n897), .B2(new_n883), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n884), .A2(new_n880), .A3(new_n883), .A4(new_n886), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n401), .B2(new_n408), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n898), .A2(G469), .A3(new_n751), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n231), .A2(new_n241), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n906), .ZN(G60));
  NAND2_X1  g732(.A1(new_n614), .A2(new_n616), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n880), .A2(new_n883), .A3(new_n886), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT54), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n925), .B2(new_n887), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT124), .B1(new_n926), .B2(new_n906), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n922), .B1(new_n909), .B2(new_n910), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n929));
  INV_X1    g743(.A(new_n906), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n919), .B1(new_n888), .B2(new_n921), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT125), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G63));
  XNOR2_X1  g751(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n897), .B2(new_n883), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n930), .B1(new_n941), .B2(new_n542), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n643), .B2(new_n941), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n314), .B2(new_n561), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n865), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n606), .B1(G898), .B2(new_n189), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NOR2_X1   g762(.A1(new_n769), .A2(new_n778), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n950));
  INV_X1    g764(.A(new_n838), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n792), .A2(new_n720), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n758), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n949), .A2(new_n189), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n480), .A2(new_n481), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n234), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n954), .B(new_n956), .C1(new_n656), .C2(new_n189), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n696), .A2(new_n951), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n682), .A2(new_n749), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n712), .C1(new_n618), .C2(new_n844), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n949), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n189), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n963), .B2(new_n956), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G72));
  NAND4_X1  g780(.A1(new_n959), .A2(new_n949), .A3(new_n865), .A4(new_n961), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  AOI22_X1  g783(.A1(new_n967), .A2(new_n969), .B1(new_n482), .B2(new_n431), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n949), .A2(new_n865), .A3(new_n950), .A4(new_n953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n447), .B1(new_n971), .B2(new_n969), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n458), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n969), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n458), .B2(new_n486), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n874), .A2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n973), .A2(new_n930), .A3(new_n977), .ZN(G57));
endmodule


