

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(KEYINPUT67), .B(n525), .ZN(n595) );
  XNOR2_X1 U550 ( .A(KEYINPUT64), .B(n521), .ZN(n642) );
  OR2_X1 U551 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n535), .ZN(n875) );
  AND2_X1 U553 ( .A1(n743), .A2(n742), .ZN(n745) );
  INV_X1 U554 ( .A(KEYINPUT32), .ZN(n744) );
  AND2_X1 U555 ( .A1(n719), .A2(n512), .ZN(n721) );
  XNOR2_X1 U556 ( .A(n690), .B(KEYINPUT31), .ZN(n691) );
  INV_X1 U557 ( .A(KEYINPUT98), .ZN(n690) );
  XNOR2_X1 U558 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U559 ( .A1(n752), .A2(n518), .ZN(n753) );
  XNOR2_X1 U560 ( .A(n588), .B(n587), .ZN(n589) );
  INV_X2 U561 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XNOR2_X1 U563 ( .A(KEYINPUT28), .B(n718), .ZN(n512) );
  NOR2_X1 U564 ( .A1(n693), .A2(n998), .ZN(n513) );
  AND2_X1 U565 ( .A1(n748), .A2(n996), .ZN(n514) );
  NOR2_X1 U566 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U567 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X2 U568 ( .A(n578), .B(n577), .ZN(G160) );
  NOR2_X1 U569 ( .A1(n802), .A2(n517), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n749), .A2(KEYINPUT33), .ZN(n516) );
  AND2_X1 U571 ( .A1(n1009), .A2(n814), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n751), .A2(KEYINPUT33), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n695), .A2(G1996), .ZN(n696) );
  XNOR2_X1 U574 ( .A(n696), .B(KEYINPUT26), .ZN(n699) );
  NOR2_X1 U575 ( .A1(G1966), .A2(n731), .ZN(n729) );
  NAND2_X1 U576 ( .A1(n730), .A2(n746), .ZN(n761) );
  INV_X1 U577 ( .A(KEYINPUT13), .ZN(n586) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  XNOR2_X1 U579 ( .A(n586), .B(KEYINPUT72), .ZN(n587) );
  OR2_X1 U580 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n646) );
  NOR2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G171) );
  INV_X1 U583 ( .A(G651), .ZN(n524) );
  NOR2_X1 U584 ( .A1(G543), .A2(n524), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n519), .Z(n520) );
  XNOR2_X2 U586 ( .A(KEYINPUT68), .B(n520), .ZN(n641) );
  NAND2_X1 U587 ( .A1(G64), .A2(n641), .ZN(n523) );
  NOR2_X1 U588 ( .A1(G651), .A2(n635), .ZN(n521) );
  NAND2_X1 U589 ( .A1(G52), .A2(n642), .ZN(n522) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n531) );
  OR2_X1 U591 ( .A1(n524), .A2(n635), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n595), .A2(G77), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT70), .ZN(n528) );
  NAND2_X1 U594 ( .A1(G90), .A2(n646), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n529), .Z(n530) );
  XOR2_X2 U597 ( .A(KEYINPUT17), .B(n532), .Z(n879) );
  NAND2_X1 U598 ( .A1(G138), .A2(n879), .ZN(n534) );
  AND2_X4 U599 ( .A1(n535), .A2(G2104), .ZN(n880) );
  NAND2_X1 U600 ( .A1(G102), .A2(n880), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n539) );
  NAND2_X1 U602 ( .A1(G126), .A2(n875), .ZN(n537) );
  AND2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U604 ( .A1(G114), .A2(n876), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(G164) );
  NAND2_X1 U607 ( .A1(n595), .A2(G78), .ZN(n541) );
  NAND2_X1 U608 ( .A1(G65), .A2(n641), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n646), .A2(G91), .ZN(n543) );
  NAND2_X1 U611 ( .A1(G53), .A2(n642), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U613 ( .A1(n545), .A2(n544), .ZN(G299) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U615 ( .A1(n875), .A2(G123), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n546), .B(KEYINPUT18), .ZN(n548) );
  NAND2_X1 U617 ( .A1(G135), .A2(n879), .ZN(n547) );
  NAND2_X1 U618 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U619 ( .A(KEYINPUT78), .B(n549), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G99), .A2(n880), .ZN(n551) );
  NAND2_X1 U621 ( .A1(G111), .A2(n876), .ZN(n550) );
  NAND2_X1 U622 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U624 ( .A(KEYINPUT79), .B(n554), .ZN(n916) );
  XNOR2_X1 U625 ( .A(G2096), .B(n916), .ZN(n555) );
  OR2_X1 U626 ( .A1(G2100), .A2(n555), .ZN(G156) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U628 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n646), .A2(G89), .ZN(n556) );
  XNOR2_X1 U630 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U631 ( .A1(G76), .A2(n595), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U633 ( .A(n559), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n564) );
  NAND2_X1 U635 ( .A1(G51), .A2(n642), .ZN(n560) );
  XNOR2_X1 U636 ( .A(n560), .B(KEYINPUT74), .ZN(n562) );
  NAND2_X1 U637 ( .A1(G63), .A2(n641), .ZN(n561) );
  NAND2_X1 U638 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U639 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U641 ( .A(n568), .B(n567), .ZN(G168) );
  XOR2_X1 U642 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U643 ( .A(KEYINPUT65), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n880), .A2(G101), .ZN(n569) );
  XOR2_X1 U645 ( .A(KEYINPUT23), .B(n569), .Z(n571) );
  NAND2_X1 U646 ( .A1(n875), .A2(G125), .ZN(n570) );
  NAND2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U648 ( .A(n572), .B(KEYINPUT66), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G137), .A2(n879), .ZN(n574) );
  NAND2_X1 U650 ( .A1(G113), .A2(n876), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n830) );
  NAND2_X1 U655 ( .A1(n830), .A2(G567), .ZN(n580) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U657 ( .A1(G56), .A2(n641), .ZN(n581) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n581), .Z(n590) );
  NAND2_X1 U659 ( .A1(G68), .A2(n595), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n583) );
  NAND2_X1 U661 ( .A1(G81), .A2(n646), .ZN(n582) );
  XNOR2_X1 U662 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n588) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G43), .A2(n642), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n998) );
  INV_X1 U667 ( .A(G860), .ZN(n606) );
  OR2_X1 U668 ( .A1(n998), .A2(n606), .ZN(G153) );
  XNOR2_X1 U669 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n646), .A2(G92), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G54), .A2(n642), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n595), .A2(G79), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G66), .A2(n641), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X2 U677 ( .A(n600), .B(KEYINPUT15), .ZN(n1003) );
  OR2_X1 U678 ( .A1(n1003), .A2(G868), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(G284) );
  INV_X1 U680 ( .A(G868), .ZN(n662) );
  NAND2_X1 U681 ( .A1(G299), .A2(n662), .ZN(n604) );
  NAND2_X1 U682 ( .A1(G868), .A2(G286), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT77), .B(n605), .Z(G297) );
  NAND2_X1 U685 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n607), .A2(n1003), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n998), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G868), .A2(n1003), .ZN(n609) );
  NOR2_X1 U690 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U692 ( .A1(n1003), .A2(G559), .ZN(n659) );
  XNOR2_X1 U693 ( .A(n998), .B(n659), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n612), .A2(G860), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n595), .A2(G80), .ZN(n614) );
  NAND2_X1 U696 ( .A1(G67), .A2(n641), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n646), .A2(G93), .ZN(n616) );
  NAND2_X1 U699 ( .A1(G55), .A2(n642), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n661) );
  XOR2_X1 U702 ( .A(n619), .B(n661), .Z(G145) );
  NAND2_X1 U703 ( .A1(n595), .A2(G75), .ZN(n621) );
  NAND2_X1 U704 ( .A1(G62), .A2(n641), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G88), .A2(n646), .ZN(n622) );
  XNOR2_X1 U707 ( .A(KEYINPUT81), .B(n622), .ZN(n623) );
  NOR2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G50), .A2(n642), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(n646), .A2(G86), .ZN(n628) );
  NAND2_X1 U713 ( .A1(G61), .A2(n641), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n595), .A2(G73), .ZN(n629) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G48), .A2(n642), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U720 ( .A1(n642), .A2(G49), .ZN(n634) );
  XNOR2_X1 U721 ( .A(n634), .B(KEYINPUT80), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U725 ( .A1(n641), .A2(n638), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G60), .A2(n641), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G47), .A2(n642), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U730 ( .A(KEYINPUT69), .B(n645), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G72), .A2(n595), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G85), .A2(n646), .ZN(n647) );
  AND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G290) );
  XNOR2_X1 U735 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n998), .B(KEYINPUT19), .ZN(n651) );
  XNOR2_X1 U737 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U738 ( .A(n661), .B(n653), .Z(n655) );
  XNOR2_X1 U739 ( .A(G299), .B(G166), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U741 ( .A(n656), .B(G305), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n657), .B(G288), .ZN(n658) );
  XNOR2_X1 U743 ( .A(n658), .B(G290), .ZN(n905) );
  XNOR2_X1 U744 ( .A(n659), .B(n905), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(G2072), .ZN(n669) );
  XNOR2_X1 U753 ( .A(KEYINPUT84), .B(n669), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n671) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U758 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U759 ( .A1(n672), .A2(G218), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G96), .A2(n673), .ZN(n834) );
  NAND2_X1 U761 ( .A1(n834), .A2(G2106), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G120), .A2(G69), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U764 ( .A1(G108), .A2(n675), .ZN(n835) );
  NAND2_X1 U765 ( .A1(n835), .A2(G567), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n836) );
  NOR2_X1 U767 ( .A1(n678), .A2(n836), .ZN(n679) );
  XNOR2_X1 U768 ( .A(n679), .B(KEYINPUT86), .ZN(n833) );
  NAND2_X1 U769 ( .A1(G36), .A2(n833), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U771 ( .A(n770), .ZN(n680) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X1 U773 ( .A1(n680), .A2(n771), .ZN(n694) );
  BUF_X2 U774 ( .A(n694), .Z(n697) );
  NAND2_X1 U775 ( .A1(n697), .A2(G8), .ZN(n681) );
  XOR2_X1 U776 ( .A(KEYINPUT91), .B(n681), .Z(n731) );
  NOR2_X1 U777 ( .A1(G2084), .A2(n697), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n729), .A2(n725), .ZN(n682) );
  NAND2_X1 U779 ( .A1(G8), .A2(n682), .ZN(n683) );
  XNOR2_X1 U780 ( .A(KEYINPUT30), .B(n683), .ZN(n684) );
  NOR2_X1 U781 ( .A1(G168), .A2(n684), .ZN(n689) );
  INV_X1 U782 ( .A(G1961), .ZN(n943) );
  NAND2_X1 U783 ( .A1(n697), .A2(n943), .ZN(n686) );
  INV_X1 U784 ( .A(n697), .ZN(n710) );
  XNOR2_X1 U785 ( .A(KEYINPUT25), .B(G2078), .ZN(n974) );
  NAND2_X1 U786 ( .A1(n710), .A2(n974), .ZN(n685) );
  NAND2_X1 U787 ( .A1(n686), .A2(n685), .ZN(n722) );
  NOR2_X1 U788 ( .A1(G171), .A2(n722), .ZN(n687) );
  XOR2_X1 U789 ( .A(KEYINPUT97), .B(n687), .Z(n688) );
  NOR2_X1 U790 ( .A1(n689), .A2(n688), .ZN(n692) );
  XNOR2_X1 U791 ( .A(n692), .B(n691), .ZN(n736) );
  INV_X1 U792 ( .A(n1003), .ZN(n693) );
  INV_X1 U793 ( .A(n694), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n697), .A2(G1341), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n706) );
  INV_X1 U796 ( .A(n706), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n513), .A2(n700), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n710), .A2(G1348), .ZN(n702) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n697), .ZN(n701) );
  NOR2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U802 ( .A(KEYINPUT94), .B(n705), .Z(n709) );
  NOR2_X1 U803 ( .A1(n998), .A2(n706), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n1003), .A2(n707), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n710), .A2(G2072), .ZN(n711) );
  XOR2_X1 U807 ( .A(KEYINPUT27), .B(n711), .Z(n713) );
  NAND2_X1 U808 ( .A1(G1956), .A2(n697), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U810 ( .A1(G299), .A2(n717), .ZN(n714) );
  XNOR2_X1 U811 ( .A(n716), .B(KEYINPUT95), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G299), .A2(n717), .ZN(n718) );
  XNOR2_X1 U813 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n721), .B(n720), .ZN(n724) );
  NAND2_X1 U815 ( .A1(G171), .A2(n722), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n738) );
  NAND2_X1 U817 ( .A1(n736), .A2(n738), .ZN(n727) );
  NAND2_X1 U818 ( .A1(G8), .A2(n725), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  INV_X1 U820 ( .A(n731), .ZN(n765) );
  INV_X1 U821 ( .A(n765), .ZN(n749) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n749), .ZN(n733) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n697), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n734), .A2(G303), .ZN(n735) );
  XOR2_X1 U826 ( .A(KEYINPUT99), .B(n735), .Z(n739) );
  AND2_X1 U827 ( .A1(n736), .A2(n739), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n743) );
  INV_X1 U829 ( .A(n739), .ZN(n740) );
  OR2_X1 U830 ( .A1(n740), .A2(G286), .ZN(n741) );
  AND2_X1 U831 ( .A1(n741), .A2(G8), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n750), .A2(n747), .ZN(n997) );
  NAND2_X1 U835 ( .A1(n761), .A2(n997), .ZN(n748) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n996) );
  NAND2_X1 U837 ( .A1(n514), .A2(n516), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n750), .A2(n765), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n753), .B(KEYINPUT100), .ZN(n754) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n993) );
  NAND2_X1 U841 ( .A1(n754), .A2(n993), .ZN(n760) );
  XOR2_X1 U842 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n755) );
  XNOR2_X1 U843 ( .A(KEYINPUT92), .B(n755), .ZN(n757) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XNOR2_X1 U845 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n758), .A2(n765), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n768) );
  INV_X1 U848 ( .A(n761), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G166), .A2(G8), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  INV_X1 U854 ( .A(n769), .ZN(n803) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n814) );
  NAND2_X1 U856 ( .A1(G140), .A2(n879), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G104), .A2(n880), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G128), .A2(n875), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G116), .A2(n876), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U863 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(KEYINPUT36), .B(n780), .ZN(n888) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NOR2_X1 U867 ( .A1(n888), .A2(n812), .ZN(n915) );
  NAND2_X1 U868 ( .A1(n814), .A2(n915), .ZN(n810) );
  NAND2_X1 U869 ( .A1(n880), .A2(G95), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT87), .B(n781), .Z(n783) );
  NAND2_X1 U871 ( .A1(n879), .A2(G131), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT88), .B(n784), .Z(n788) );
  NAND2_X1 U874 ( .A1(G119), .A2(n875), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G107), .A2(n876), .ZN(n785) );
  AND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n893) );
  AND2_X1 U878 ( .A1(n893), .A2(G1991), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G129), .A2(n875), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G117), .A2(n876), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n880), .A2(G105), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT89), .B(n794), .Z(n796) );
  NAND2_X1 U886 ( .A1(n879), .A2(G141), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n894) );
  AND2_X1 U888 ( .A1(n894), .A2(G1996), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n925) );
  INV_X1 U890 ( .A(n814), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n925), .A2(n799), .ZN(n806) );
  INV_X1 U892 ( .A(n806), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n810), .A2(n800), .ZN(n801) );
  XNOR2_X1 U894 ( .A(KEYINPUT90), .B(n801), .ZN(n802) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n1009) );
  NAND2_X1 U896 ( .A1(n803), .A2(n515), .ZN(n817) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n894), .ZN(n933) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n893), .ZN(n914) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n804) );
  XOR2_X1 U900 ( .A(n804), .B(KEYINPUT101), .Z(n805) );
  NOR2_X1 U901 ( .A1(n914), .A2(n805), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U903 ( .A1(n933), .A2(n808), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n888), .A2(n812), .ZN(n924) );
  NAND2_X1 U907 ( .A1(n813), .A2(n924), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  XNOR2_X1 U911 ( .A(G2427), .B(G2451), .ZN(n828) );
  XOR2_X1 U912 ( .A(G2430), .B(G2443), .Z(n820) );
  XNOR2_X1 U913 ( .A(G2435), .B(KEYINPUT102), .ZN(n819) );
  XNOR2_X1 U914 ( .A(n820), .B(n819), .ZN(n824) );
  XOR2_X1 U915 ( .A(G2438), .B(G2454), .Z(n822) );
  XNOR2_X1 U916 ( .A(G1341), .B(G1348), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U918 ( .A(n824), .B(n823), .Z(n826) );
  XNOR2_X1 U919 ( .A(KEYINPUT103), .B(G2446), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(G14), .ZN(n908) );
  XOR2_X1 U923 ( .A(KEYINPUT104), .B(n908), .Z(G401) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  XOR2_X1 U930 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  NOR2_X1 U935 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n836), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT109), .B(G1966), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U941 ( .A(n839), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1971), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U944 ( .A(G1976), .B(G1981), .Z(n843) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT110), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n849) );
  XNOR2_X1 U951 ( .A(G2678), .B(KEYINPUT43), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U953 ( .A(KEYINPUT42), .B(G2090), .Z(n851) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U956 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U957 ( .A(G2096), .B(G2100), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U959 ( .A(G2084), .B(G2078), .Z(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(G227) );
  NAND2_X1 U961 ( .A1(G124), .A2(n875), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n880), .A2(G100), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G136), .A2(n879), .ZN(n862) );
  NAND2_X1 U966 ( .A1(G112), .A2(n876), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U968 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U969 ( .A1(n880), .A2(G103), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n865), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G139), .A2(n879), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U973 ( .A(KEYINPUT113), .B(n868), .Z(n874) );
  NAND2_X1 U974 ( .A1(n876), .A2(G115), .ZN(n869) );
  XNOR2_X1 U975 ( .A(n869), .B(KEYINPUT114), .ZN(n871) );
  NAND2_X1 U976 ( .A1(G127), .A2(n875), .ZN(n870) );
  NAND2_X1 U977 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n918) );
  NAND2_X1 U980 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n918), .B(n886), .ZN(n898) );
  XOR2_X1 U989 ( .A(G164), .B(G162), .Z(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n890) );
  XNOR2_X1 U992 ( .A(KEYINPUT115), .B(KEYINPUT111), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(n892), .B(n891), .Z(n896) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n916), .B(G160), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(G286), .B(KEYINPUT116), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G171), .B(n1003), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT117), .B(n907), .Z(G397) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n908), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n939) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n931) );
  XNOR2_X1 U1018 ( .A(G2072), .B(n918), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT119), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G2078), .B(G164), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n922), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n923), .B(KEYINPUT120), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT118), .B(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n935), .Z(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n939), .B(n938), .ZN(n941) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(G29), .ZN(n991) );
  XNOR2_X1 U1038 ( .A(G5), .B(n943), .ZN(n956) );
  XNOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(G4), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G20), .B(G1956), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT127), .B(G1981), .Z(n949) );
  XNOR2_X1 U1046 ( .A(G6), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT60), .B(n952), .Z(n954) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G23), .B(G1976), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1059 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1060 ( .A1(G16), .A2(n965), .ZN(n989) );
  XOR2_X1 U1061 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n984) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G35), .ZN(n979) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G32), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(G33), .B(G2072), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n973) );
  XOR2_X1 U1066 ( .A(G2067), .B(G26), .Z(n968) );
  NAND2_X1 U1067 ( .A1(n968), .A2(G28), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G25), .B(G1991), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(KEYINPUT122), .B(n969), .ZN(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1072 ( .A(G27), .B(n974), .Z(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n977), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n980), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n984), .B(n983), .ZN(n985) );
  OR2_X1 U1080 ( .A1(G29), .A2(n985), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n986), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n987), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n1018) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT125), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT56), .ZN(n1016) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT57), .B(n995), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G171), .B(G1961), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(n1003), .B(G1348), .Z(n1005) );
  XNOR2_X1 U1096 ( .A(G299), .B(G1956), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1014), .B(KEYINPUT126), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

