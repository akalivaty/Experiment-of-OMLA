//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n202), .B2(G1gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n203), .B(new_n205), .C1(new_n208), .C2(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT90), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT90), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(G64gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(G64gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT93), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  INV_X1    g022(.A(G71gat), .ZN(new_n224));
  INV_X1    g023(.A(G78gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT9), .B1(new_n217), .B2(new_n220), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n223), .A3(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n215), .B1(KEYINPUT21), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G155gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G231gat), .ZN(new_n240));
  INV_X1    g039(.A(G233gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(G231gat), .B(G233gat), .C1(new_n233), .C2(new_n238), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n237), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n236), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n248), .A2(new_n244), .A3(new_n235), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n234), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n235), .B1(new_n248), .B2(new_n244), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n246), .A3(new_n236), .ZN(new_n252));
  INV_X1    g051(.A(new_n234), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G183gat), .B(G211gat), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G190gat), .B(G218gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G99gat), .B(G106gat), .ZN(new_n262));
  INV_X1    g061(.A(G92gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT95), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT95), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G92gat), .ZN(new_n266));
  INV_X1    g065(.A(G85gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G99gat), .ZN(new_n269));
  INV_X1    g068(.A(G106gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT8), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT96), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT96), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G85gat), .A2(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT7), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n262), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n268), .A2(new_n274), .A3(new_n271), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n268), .B2(new_n271), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n262), .B(new_n278), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT17), .ZN(new_n285));
  NAND2_X1  g084(.A1(G29gat), .A2(G36gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT15), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G43gat), .B(G50gat), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT15), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n290), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT15), .A3(new_n293), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n285), .B1(new_n299), .B2(KEYINPUT88), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n298), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT17), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n284), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n307));
  INV_X1    g106(.A(new_n262), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n282), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n310), .B2(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n261), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT17), .B1(new_n301), .B2(new_n302), .ZN(new_n314));
  AOI211_X1 g113(.A(KEYINPUT88), .B(new_n285), .C1(new_n296), .C2(new_n298), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n261), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n322));
  XNOR2_X1  g121(.A(G134gat), .B(G162gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n312), .B(new_n318), .C1(new_n320), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G230gat), .A2(G233gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n330), .B(KEYINPUT98), .Z(new_n331));
  OAI21_X1  g130(.A(new_n232), .B1(new_n279), .B2(new_n283), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n309), .A2(new_n233), .A3(new_n282), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n284), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n331), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G120gat), .B(G148gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G176gat), .B(G204gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n344), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n260), .A2(new_n329), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G78gat), .B(G106gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT78), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT31), .B(G50gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT79), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n358), .B(new_n364), .C1(new_n361), .C2(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  INV_X1    g169(.A(G148gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G155gat), .B(G162gat), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G155gat), .B(G162gat), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n372), .A2(new_n381), .A3(new_n373), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT73), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT73), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n357), .B1(new_n369), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n367), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n357), .B(new_n385), .C1(new_n368), .C2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n356), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n369), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n355), .B1(new_n388), .B2(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n354), .B1(new_n401), .B2(KEYINPUT81), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(G22gat), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n408));
  INV_X1    g207(.A(new_n384), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT73), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n392), .A3(new_n391), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(new_n356), .B1(new_n399), .B2(new_n398), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n414), .B2(new_n403), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n402), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(G22gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n403), .A3(new_n406), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n414), .A2(new_n403), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n354), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT25), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT66), .B(G190gat), .ZN(new_n424));
  INV_X1    g223(.A(G183gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n423), .A3(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT24), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT64), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT64), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(G169gat), .A3(G176gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(G169gat), .A2(G176gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT23), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT65), .B1(new_n433), .B2(new_n435), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n422), .B1(new_n431), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(G183gat), .B2(G190gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n439), .B(KEYINPUT23), .Z(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(new_n422), .A3(new_n436), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n439), .A2(KEYINPUT26), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT26), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G169gat), .B2(G176gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n450), .A2(new_n436), .B1(G183gat), .B2(G190gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT27), .B(G183gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n452), .A3(KEYINPUT28), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT28), .B1(new_n424), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT72), .B1(new_n443), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n453), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n433), .A2(new_n435), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n440), .A2(new_n461), .A3(KEYINPUT25), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n460), .A2(new_n451), .B1(new_n462), .B2(new_n444), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n428), .A2(new_n430), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n426), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(KEYINPUT65), .ZN(new_n466));
  INV_X1    g265(.A(new_n441), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n445), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT25), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT29), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n463), .A2(new_n469), .A3(new_n472), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n390), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n458), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n469), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n481), .A2(new_n472), .B1(new_n473), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n476), .B(new_n480), .C1(new_n483), .C2(new_n390), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n476), .B(new_n485), .C1(new_n483), .C2(new_n390), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n479), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n474), .A2(new_n389), .A3(new_n475), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT37), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n443), .A2(new_n457), .A3(KEYINPUT72), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n470), .B1(new_n463), .B2(new_n469), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n472), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n482), .A2(new_n473), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n389), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n488), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n484), .B1(new_n487), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n390), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n474), .A2(new_n390), .A3(new_n475), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT37), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n479), .A3(new_n486), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(KEYINPUT38), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  XOR2_X1   g302(.A(G1gat), .B(G29gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT0), .ZN(new_n505));
  XNOR2_X1  g304(.A(G57gat), .B(G85gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT1), .ZN(new_n509));
  INV_X1    g308(.A(G113gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(G120gat), .ZN(new_n511));
  INV_X1    g310(.A(G120gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(G113gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n515), .A2(new_n509), .B1(G127gat), .B2(G134gat), .ZN(new_n516));
  OR2_X1    g315(.A1(G127gat), .A2(G134gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n514), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n395), .A2(new_n520), .A3(new_n397), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n411), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G225gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n508), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n525), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n521), .B2(new_n522), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT77), .B1(new_n530), .B2(new_n508), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT4), .B1(new_n520), .B2(new_n385), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n522), .A2(new_n534), .A3(KEYINPUT4), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n411), .A2(new_n536), .A3(new_n519), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n395), .A2(KEYINPUT3), .A3(new_n397), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT3), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n519), .B1(new_n411), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n525), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n531), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n532), .A2(new_n537), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n547), .A2(KEYINPUT5), .A3(new_n525), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n503), .B(new_n507), .C1(new_n544), .C2(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n526), .A2(new_n527), .B1(new_n538), .B2(new_n542), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n551), .B2(new_n531), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT6), .B1(new_n552), .B2(new_n507), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n544), .A2(new_n549), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n507), .B(KEYINPUT82), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n550), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n421), .B1(new_n502), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n484), .A2(KEYINPUT30), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n479), .B1(new_n498), .B2(new_n499), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT30), .A3(new_n484), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n539), .A2(new_n541), .B1(new_n532), .B2(new_n537), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n566), .A2(KEYINPUT39), .A3(new_n529), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n567), .B2(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n525), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT83), .B(new_n555), .C1(new_n569), .C2(KEYINPUT39), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n566), .A2(new_n529), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT39), .B1(new_n523), .B2(new_n525), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT40), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n577), .B(new_n574), .C1(new_n568), .C2(new_n570), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT84), .B1(new_n564), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT84), .ZN(new_n581));
  NOR4_X1   g380(.A1(new_n563), .A2(new_n576), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n559), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n507), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n503), .B1(new_n554), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n552), .A2(new_n507), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n560), .A2(new_n562), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n520), .B1(new_n443), .B2(new_n457), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n463), .A2(new_n469), .A3(new_n519), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G227gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n241), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT32), .ZN(new_n598));
  XOR2_X1   g397(.A(G15gat), .B(G43gat), .Z(new_n599));
  XNOR2_X1  g398(.A(G71gat), .B(G99gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n601), .B2(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(KEYINPUT69), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT69), .ZN(new_n604));
  INV_X1    g403(.A(new_n596), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n592), .B2(new_n593), .ZN(new_n606));
  INV_X1    g405(.A(new_n602), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n597), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n601), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n593), .A3(new_n605), .ZN(new_n614));
  OR3_X1    g413(.A1(new_n614), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT70), .B1(new_n614), .B2(KEYINPUT34), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(KEYINPUT34), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n613), .A2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n591), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(KEYINPUT36), .A3(new_n619), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n590), .A2(new_n421), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT86), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n560), .A2(new_n562), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n558), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n552), .A2(new_n555), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n585), .B1(new_n586), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(KEYINPUT86), .A3(new_n589), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n416), .A2(new_n420), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n603), .A2(new_n608), .B1(new_n611), .B2(new_n601), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n618), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n588), .A2(new_n589), .A3(new_n635), .A4(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT35), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT92), .ZN(new_n643));
  XNOR2_X1  g442(.A(G113gat), .B(G141gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT11), .ZN(new_n645));
  INV_X1    g444(.A(G169gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G197gat), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n648), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n212), .B1(new_n314), .B2(new_n315), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n213), .A2(new_n301), .A3(new_n215), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(KEYINPUT91), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n654), .B(KEYINPUT13), .Z(new_n659));
  INV_X1    g458(.A(new_n655), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n301), .B1(new_n213), .B2(new_n215), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n657), .B1(new_n656), .B2(KEYINPUT91), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n652), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(KEYINPUT91), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT18), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(new_n651), .A3(new_n658), .A4(new_n662), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n642), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n583), .A2(new_n625), .B1(new_n638), .B2(new_n640), .ZN(new_n671));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT92), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n350), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n588), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g476(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n204), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(new_n628), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G8gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(G8gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n674), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n589), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n681), .B(new_n682), .C1(KEYINPUT42), .C2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(new_n635), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n683), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n622), .A2(new_n624), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT100), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n622), .A2(new_n624), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n687), .A2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n674), .A2(new_n421), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n260), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n328), .A3(new_n349), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n588), .A2(G29gat), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n701), .B(new_n702), .C1(new_n670), .C2(new_n673), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n671), .B2(new_n329), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n554), .A2(new_n584), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n553), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n628), .B1(new_n585), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n690), .B1(new_n710), .B2(new_n633), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n576), .A2(new_n578), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n581), .B1(new_n712), .B2(new_n563), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n564), .A2(new_n579), .A3(KEYINPUT84), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n715), .B2(new_n559), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n553), .A2(new_n557), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n718), .A2(new_n585), .B1(new_n562), .B2(new_n560), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(KEYINPUT86), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n720), .A2(new_n629), .B1(KEYINPUT35), .B2(new_n639), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n328), .C1(new_n716), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n260), .B(KEYINPUT103), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n669), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n668), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n723), .A2(new_n348), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n722), .A3(new_n675), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G29gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n704), .B(new_n705), .C1(new_n730), .C2(new_n732), .ZN(G1328gat));
  NAND3_X1  g532(.A1(new_n707), .A2(new_n722), .A3(new_n728), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n734), .B2(new_n589), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n701), .B1(new_n670), .B2(new_n673), .ZN(new_n736));
  INV_X1    g535(.A(G36gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n628), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT46), .B1(new_n736), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(G1329gat));
  OAI21_X1  g541(.A(G43gat), .B1(new_n734), .B2(new_n690), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n686), .A2(G43gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n745), .A3(KEYINPUT47), .ZN(new_n746));
  INV_X1    g545(.A(new_n693), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n707), .A2(new_n722), .A3(new_n747), .A4(new_n728), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n736), .A2(new_n744), .B1(new_n748), .B2(G43gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(KEYINPUT47), .B2(new_n749), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n421), .A2(G50gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n707), .A2(new_n722), .A3(new_n728), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n736), .A2(new_n421), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n753), .B(new_n758), .C1(new_n759), .C2(G50gat), .ZN(new_n760));
  AOI21_X1  g559(.A(G50gat), .B1(new_n736), .B2(new_n421), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n751), .B(new_n752), .C1(new_n761), .C2(new_n757), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n760), .A2(new_n762), .ZN(G1331gat));
  AND2_X1   g562(.A1(new_n725), .A2(new_n726), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n699), .A2(new_n764), .A3(new_n328), .A4(new_n349), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n642), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n588), .B(KEYINPUT106), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT107), .B(G57gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1332gat));
  INV_X1    g570(.A(new_n766), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n628), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n774), .B2(new_n773), .ZN(G1333gat));
  OAI21_X1  g576(.A(new_n224), .B1(new_n766), .B2(new_n686), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n747), .A2(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n633), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n225), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n764), .A2(new_n260), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n348), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n707), .A2(new_n722), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n707), .A2(new_n722), .A3(KEYINPUT108), .A4(new_n786), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n675), .A3(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n328), .B(new_n784), .C1(new_n716), .C2(new_n721), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n642), .A2(KEYINPUT51), .A3(new_n328), .A4(new_n784), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n675), .A2(new_n267), .A3(new_n348), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n791), .A2(new_n267), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  NAND4_X1  g598(.A1(new_n707), .A2(new_n722), .A3(new_n628), .A4(new_n786), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n264), .A2(new_n266), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n349), .A2(G92gat), .A3(new_n589), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n796), .A2(KEYINPUT109), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT109), .B1(new_n796), .B2(new_n803), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n628), .A3(new_n790), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(new_n801), .B1(new_n796), .B2(new_n803), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n747), .A3(new_n790), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n789), .A2(new_n813), .A3(new_n747), .A4(new_n790), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(G99gat), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n269), .A3(new_n635), .A4(new_n348), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1338gat));
  NOR3_X1   g616(.A1(new_n349), .A2(new_n633), .A3(G106gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT111), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n796), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT113), .B1(new_n787), .B2(new_n633), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n633), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n789), .A2(new_n421), .A3(new_n790), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n819), .B(KEYINPUT112), .Z(new_n826));
  AOI22_X1  g625(.A1(new_n825), .A2(G106gat), .B1(new_n796), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  NOR2_X1   g628(.A1(new_n350), .A2(new_n764), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n335), .A2(new_n336), .ZN(new_n833));
  INV_X1    g632(.A(new_n331), .ZN(new_n834));
  XOR2_X1   g633(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n344), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n335), .A2(new_n336), .A3(new_n331), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n335), .A2(new_n336), .A3(new_n840), .A4(new_n331), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n337), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n832), .B1(new_n845), .B2(KEYINPUT55), .ZN(new_n846));
  INV_X1    g645(.A(new_n661), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n655), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n848), .A2(new_n659), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n648), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n328), .A2(new_n668), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n842), .A2(new_n844), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT116), .B(new_n855), .C1(new_n856), .C2(new_n837), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n345), .B1(new_n845), .B2(KEYINPUT55), .ZN(new_n858));
  AND4_X1   g657(.A1(new_n846), .A2(new_n854), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n348), .A2(new_n668), .A3(new_n853), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n846), .A3(new_n858), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n727), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n329), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n831), .B1(new_n863), .B2(new_n723), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n421), .A2(new_n686), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n675), .A3(new_n589), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n510), .A3(new_n672), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n865), .A3(new_n767), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT118), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n864), .A2(new_n871), .A3(new_n865), .A4(new_n767), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n589), .A3(new_n764), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n510), .ZN(G1340gat));
  NOR3_X1   g674(.A1(new_n867), .A2(new_n512), .A3(new_n349), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n873), .A2(new_n589), .A3(new_n348), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n512), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n723), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n867), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n628), .B(new_n699), .C1(new_n870), .C2(new_n872), .ZN(new_n882));
  AOI21_X1  g681(.A(G127gat), .B1(new_n882), .B2(KEYINPUT119), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n873), .A2(new_n589), .A3(new_n260), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n881), .B1(new_n883), .B2(new_n886), .ZN(G1342gat));
  OAI21_X1  g686(.A(G134gat), .B1(new_n867), .B2(new_n329), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n628), .A2(G134gat), .A3(new_n329), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n873), .A2(KEYINPUT56), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT56), .B1(new_n873), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n747), .A2(new_n768), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n864), .A3(new_n589), .A4(new_n421), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n672), .A2(G141gat), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT58), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n688), .A2(new_n588), .A3(new_n628), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n864), .B2(new_n421), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n633), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n842), .A2(new_n844), .ZN(new_n904));
  INV_X1    g703(.A(new_n837), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(KEYINPUT55), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n346), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n845), .A2(KEYINPUT55), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n855), .B1(new_n856), .B2(new_n837), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n858), .A2(new_n910), .A3(KEYINPUT120), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n669), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n328), .B1(new_n912), .B2(new_n860), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n699), .B1(new_n913), .B2(new_n859), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n902), .B1(new_n914), .B2(new_n831), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n669), .B(new_n898), .C1(new_n899), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G141gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n897), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n898), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n862), .A2(new_n329), .ZN(new_n923));
  INV_X1    g722(.A(new_n859), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n830), .B1(new_n925), .B2(new_n880), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n900), .B1(new_n926), .B2(new_n633), .ZN(new_n927));
  INV_X1    g726(.A(new_n915), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n370), .B1(new_n929), .B2(new_n764), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n895), .A2(new_n931), .A3(new_n896), .ZN(new_n932));
  INV_X1    g731(.A(new_n896), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT121), .B1(new_n894), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT58), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n936), .ZN(G1344gat));
  NAND3_X1  g736(.A1(new_n895), .A2(new_n371), .A3(new_n348), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n348), .B(new_n898), .C1(new_n899), .C2(new_n915), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n371), .A2(KEYINPUT59), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(KEYINPUT123), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n914), .B1(new_n669), .B2(new_n350), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n947), .B2(new_n421), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n926), .A2(new_n900), .A3(new_n633), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n348), .B(new_n898), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n938), .B1(new_n945), .B2(new_n951), .ZN(G1345gat));
  INV_X1    g751(.A(new_n929), .ZN(new_n953));
  OAI21_X1  g752(.A(G155gat), .B1(new_n953), .B2(new_n880), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n260), .A2(new_n376), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n894), .B2(new_n955), .ZN(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n953), .B2(new_n329), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n864), .A2(new_n421), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n893), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n589), .A2(new_n377), .A3(new_n328), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n675), .A2(new_n589), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n866), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n764), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n767), .A2(new_n589), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n864), .A2(new_n865), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n864), .A2(KEYINPUT124), .A3(new_n865), .A4(new_n966), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n672), .A2(new_n646), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  INV_X1    g772(.A(G176gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n964), .A2(new_n974), .A3(new_n348), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n971), .A2(new_n348), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(G1349gat));
  NAND3_X1  g776(.A1(new_n969), .A2(new_n723), .A3(new_n970), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G183gat), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n260), .A2(new_n452), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n864), .A2(new_n865), .A3(new_n962), .A4(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT125), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT60), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT60), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n979), .A2(new_n985), .A3(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1350gat));
  NAND3_X1  g786(.A1(new_n964), .A2(new_n424), .A3(new_n328), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n328), .A3(new_n970), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n989), .A2(new_n990), .A3(G190gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n989), .B2(G190gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1351gat));
  OR2_X1    g792(.A1(new_n948), .A2(new_n949), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n693), .A2(new_n966), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n994), .A2(new_n669), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G197gat), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n693), .A2(new_n962), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n727), .A2(G197gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n958), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n997), .A2(new_n1001), .ZN(G1352gat));
  OAI211_X1 g801(.A(new_n348), .B(new_n995), .C1(new_n948), .C2(new_n949), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G204gat), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n958), .A2(new_n998), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n349), .A2(G204gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n958), .A2(new_n998), .A3(new_n1006), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1007), .A2(KEYINPUT62), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT62), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(G1353gat));
  INV_X1    g812(.A(new_n1005), .ZN(new_n1014));
  OR3_X1    g813(.A1(new_n1014), .A2(G211gat), .A3(new_n699), .ZN(new_n1015));
  OAI211_X1 g814(.A(new_n260), .B(new_n995), .C1(new_n948), .C2(new_n949), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1016), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1016), .B2(G211gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(G1354gat));
  NAND3_X1  g818(.A1(new_n994), .A2(new_n328), .A3(new_n995), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(G218gat), .ZN(new_n1021));
  OR3_X1    g820(.A1(new_n1014), .A2(G218gat), .A3(new_n329), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(new_n1022), .ZN(G1355gat));
endmodule


