

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n425) );
  XNOR2_X1 U325 ( .A(n426), .B(n425), .ZN(n427) );
  INV_X1 U326 ( .A(n400), .ZN(n358) );
  XNOR2_X1 U327 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U328 ( .A(n361), .B(n360), .ZN(n420) );
  XNOR2_X1 U329 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n463) );
  NOR2_X1 U330 ( .A1(n540), .A2(n454), .ZN(n572) );
  XNOR2_X1 U331 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U332 ( .A(n455), .B(G176GAT), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n359) );
  XOR2_X1 U335 ( .A(G127GAT), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n442) );
  XOR2_X1 U338 ( .A(n359), .B(n442), .Z(n295) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U341 ( .A(n296), .B(G183GAT), .Z(n300) );
  XOR2_X1 U342 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n336) );
  XNOR2_X1 U345 ( .A(n336), .B(KEYINPUT64), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT84), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G99GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U350 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT88), .Z(n306) );
  XNOR2_X1 U352 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U354 ( .A(G176GAT), .B(KEYINPUT20), .Z(n308) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G15GAT), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n540) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(G78GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n313), .B(G148GAT), .ZN(n344) );
  XOR2_X1 U361 ( .A(G204GAT), .B(n344), .Z(n315) );
  XOR2_X1 U362 ( .A(G141GAT), .B(G22GAT), .Z(n369) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(n369), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n331) );
  XOR2_X1 U368 ( .A(n331), .B(KEYINPUT91), .Z(n319) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U371 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U372 ( .A(KEYINPUT89), .B(G162GAT), .Z(n323) );
  XNOR2_X1 U373 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT3), .B(n324), .Z(n451) );
  XOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n326) );
  XNOR2_X1 U377 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n451), .B(n327), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n477) );
  XOR2_X1 U381 ( .A(G183GAT), .B(KEYINPUT76), .Z(n388) );
  XOR2_X1 U382 ( .A(G190GAT), .B(KEYINPUT75), .Z(n399) );
  XOR2_X1 U383 ( .A(n388), .B(n399), .Z(n333) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(G36GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n330), .B(G8GAT), .ZN(n366) );
  XNOR2_X1 U386 ( .A(n366), .B(n331), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n341) );
  XOR2_X1 U388 ( .A(G64GAT), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n355) );
  XOR2_X1 U391 ( .A(KEYINPUT96), .B(n336), .Z(n338) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(n355), .B(n339), .Z(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n528) );
  XNOR2_X1 U396 ( .A(n344), .B(KEYINPUT72), .ZN(n342) );
  AND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  NAND2_X1 U398 ( .A1(n342), .A2(n345), .ZN(n349) );
  INV_X1 U399 ( .A(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n347) );
  INV_X1 U401 ( .A(n345), .ZN(n346) );
  NAND2_X1 U402 ( .A1(n347), .A2(n346), .ZN(n348) );
  NAND2_X1 U403 ( .A1(n349), .A2(n348), .ZN(n353) );
  XOR2_X1 U404 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n351) );
  XNOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT71), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U408 ( .A(G57GAT), .B(KEYINPUT70), .Z(n354) );
  XOR2_X1 U409 ( .A(KEYINPUT13), .B(n354), .Z(n397) );
  XOR2_X1 U410 ( .A(n355), .B(n397), .Z(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n361) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G85GAT), .ZN(n400) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n363) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U416 ( .A(n364), .B(KEYINPUT30), .Z(n368) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G1GAT), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(KEYINPUT68), .ZN(n396) );
  XNOR2_X1 U419 ( .A(n366), .B(n396), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U421 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U422 ( .A(G113GAT), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT8), .B(G50GAT), .Z(n374) );
  XNOR2_X1 U425 ( .A(G43GAT), .B(G29GAT), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U427 ( .A(KEYINPUT7), .B(n375), .ZN(n413) );
  XNOR2_X1 U428 ( .A(n376), .B(n413), .ZN(n575) );
  XNOR2_X1 U429 ( .A(KEYINPUT69), .B(n575), .ZN(n566) );
  XOR2_X1 U430 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n417) );
  XOR2_X1 U431 ( .A(G64GAT), .B(G155GAT), .Z(n378) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G22GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n380) );
  XNOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U437 ( .A(n382), .B(n381), .Z(n394) );
  XOR2_X1 U438 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n384) );
  XNOR2_X1 U439 ( .A(KEYINPUT77), .B(KEYINPUT79), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U441 ( .A(G78GAT), .B(G211GAT), .Z(n386) );
  XNOR2_X1 U442 ( .A(G71GAT), .B(G127GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U444 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n585) );
  INV_X1 U451 ( .A(n585), .ZN(n569) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U453 ( .A(G162GAT), .B(G218GAT), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U455 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n404) );
  XNOR2_X1 U456 ( .A(G36GAT), .B(G92GAT), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U458 ( .A(n406), .B(n405), .Z(n408) );
  XNOR2_X1 U459 ( .A(G134GAT), .B(G106GAT), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U461 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n410) );
  NAND2_X1 U462 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U464 ( .A(n412), .B(n411), .Z(n415) );
  XOR2_X1 U465 ( .A(n413), .B(KEYINPUT66), .Z(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n571) );
  XNOR2_X1 U467 ( .A(KEYINPUT36), .B(n571), .ZN(n495) );
  NAND2_X1 U468 ( .A1(n569), .A2(n495), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n418) );
  NOR2_X1 U470 ( .A1(n566), .A2(n418), .ZN(n419) );
  NAND2_X1 U471 ( .A1(n420), .A2(n419), .ZN(n428) );
  XOR2_X1 U472 ( .A(KEYINPUT41), .B(n420), .Z(n557) );
  NOR2_X1 U473 ( .A1(n575), .A2(n557), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n421), .B(KEYINPUT46), .ZN(n422) );
  NOR2_X1 U475 ( .A1(n422), .A2(n569), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT113), .ZN(n424) );
  NOR2_X1 U477 ( .A1(n424), .A2(n571), .ZN(n426) );
  NAND2_X1 U478 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U479 ( .A(KEYINPUT48), .B(n429), .ZN(n552) );
  NAND2_X1 U480 ( .A1(n528), .A2(n552), .ZN(n432) );
  XNOR2_X1 U481 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n430), .B(KEYINPUT54), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n460) );
  XOR2_X1 U484 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n434) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U487 ( .A(KEYINPUT94), .B(n435), .ZN(n449) );
  XOR2_X1 U488 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n437) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(KEYINPUT1), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U491 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n439) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(G57GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n447) );
  XOR2_X1 U495 ( .A(G85GAT), .B(G148GAT), .Z(n444) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(G120GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n501) );
  NAND2_X1 U502 ( .A1(n460), .A2(n501), .ZN(n452) );
  NOR2_X1 U503 ( .A1(n477), .A2(n452), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n557), .B(KEYINPUT107), .ZN(n542) );
  NAND2_X1 U506 ( .A1(n572), .A2(n542), .ZN(n457) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n455) );
  INV_X1 U508 ( .A(n501), .ZN(n553) );
  NAND2_X1 U509 ( .A1(n477), .A2(n540), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n458), .B(KEYINPUT26), .ZN(n470) );
  NOR2_X1 U511 ( .A1(n553), .A2(n470), .ZN(n459) );
  AND2_X1 U512 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT121), .ZN(n584) );
  INV_X1 U514 ( .A(n584), .ZN(n462) );
  NAND2_X1 U515 ( .A1(n462), .A2(n495), .ZN(n464) );
  XOR2_X1 U516 ( .A(G218GAT), .B(KEYINPUT126), .Z(n465) );
  XNOR2_X1 U517 ( .A(n466), .B(n465), .ZN(G1355GAT) );
  NAND2_X1 U518 ( .A1(n566), .A2(n420), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT73), .B(n467), .Z(n498) );
  XOR2_X1 U520 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n469) );
  INV_X1 U521 ( .A(n571), .ZN(n564) );
  NAND2_X1 U522 ( .A1(n569), .A2(n564), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n469), .B(n468), .ZN(n483) );
  XOR2_X1 U524 ( .A(KEYINPUT27), .B(n528), .Z(n478) );
  NOR2_X1 U525 ( .A1(n470), .A2(n478), .ZN(n555) );
  INV_X1 U526 ( .A(n528), .ZN(n505) );
  NOR2_X1 U527 ( .A1(n540), .A2(n505), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n477), .A2(n471), .ZN(n472) );
  XOR2_X1 U529 ( .A(n472), .B(KEYINPUT25), .Z(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT98), .B(n473), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n555), .A2(n474), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(n475), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n476), .A2(n501), .ZN(n482) );
  XOR2_X1 U534 ( .A(n477), .B(KEYINPUT28), .Z(n511) );
  INV_X1 U535 ( .A(n511), .ZN(n532) );
  OR2_X1 U536 ( .A1(n478), .A2(n532), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n501), .A2(n479), .ZN(n538) );
  NAND2_X1 U538 ( .A1(n540), .A2(n538), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT97), .B(n480), .Z(n481) );
  NAND2_X1 U540 ( .A1(n482), .A2(n481), .ZN(n494) );
  NAND2_X1 U541 ( .A1(n483), .A2(n494), .ZN(n513) );
  NOR2_X1 U542 ( .A1(n498), .A2(n513), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n491), .A2(n553), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n528), .A2(n491), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(KEYINPUT100), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n489) );
  INV_X1 U550 ( .A(n540), .ZN(n530) );
  NAND2_X1 U551 ( .A1(n491), .A2(n530), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NAND2_X1 U554 ( .A1(n532), .A2(n491), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n494), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n569), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n497), .ZN(n526) );
  NOR2_X1 U560 ( .A1(n526), .A2(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n510) );
  NOR2_X1 U563 ( .A1(n510), .A2(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n505), .A2(n510), .ZN(n506) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n508) );
  NOR2_X1 U570 ( .A1(n540), .A2(n510), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  XOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT106), .Z(n515) );
  NAND2_X1 U576 ( .A1(n575), .A2(n542), .ZN(n525) );
  NOR2_X1 U577 ( .A1(n525), .A2(n513), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n553), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n528), .A2(n521), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT109), .Z(n520) );
  NAND2_X1 U585 ( .A1(n521), .A2(n530), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n532), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n533), .A2(n553), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n528), .A2(n533), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n533), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n537) );
  XOR2_X1 U599 ( .A(G106GAT), .B(KEYINPUT111), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n552), .A2(n538), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n566), .A2(n549), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U608 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n547) );
  NAND2_X1 U612 ( .A1(n549), .A2(n569), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n571), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  AND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n575), .A2(n563), .ZN(n556) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  NOR2_X1 U622 ( .A1(n563), .A2(n557), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n585), .A2(n563), .ZN(n562) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n572), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n572), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n574), .ZN(G1351GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n584), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n577) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n584), .A2(n420), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(G1354GAT) );
endmodule

