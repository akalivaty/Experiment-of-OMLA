

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  NOR2_X1 U326 ( .A1(n572), .A2(n463), .ZN(n535) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U328 ( .A(n419), .B(n418), .ZN(n427) );
  XOR2_X1 U329 ( .A(n415), .B(n414), .Z(n294) );
  XNOR2_X1 U330 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n295) );
  XOR2_X1 U331 ( .A(n404), .B(KEYINPUT85), .Z(n296) );
  XOR2_X1 U332 ( .A(KEYINPUT106), .B(n500), .Z(n297) );
  XNOR2_X1 U333 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n403) );
  XNOR2_X1 U334 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U335 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U336 ( .A(n394), .B(n393), .ZN(n532) );
  XNOR2_X1 U337 ( .A(n416), .B(n294), .ZN(n419) );
  INV_X1 U338 ( .A(KEYINPUT37), .ZN(n492) );
  XNOR2_X1 U339 ( .A(n361), .B(n360), .ZN(n566) );
  XNOR2_X1 U340 ( .A(n493), .B(n492), .ZN(n522) );
  XOR2_X1 U341 ( .A(n468), .B(KEYINPUT28), .Z(n528) );
  XNOR2_X1 U342 ( .A(KEYINPUT92), .B(n473), .ZN(n572) );
  XNOR2_X1 U343 ( .A(n455), .B(n295), .ZN(n456) );
  XNOR2_X1 U344 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n299) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n300), .B(KEYINPUT18), .Z(n302) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n406) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n303), .B(G127GAT), .ZN(n442) );
  XOR2_X1 U353 ( .A(n442), .B(G176GAT), .Z(n305) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n406), .B(n306), .ZN(n311) );
  XOR2_X1 U357 ( .A(G43GAT), .B(G134GAT), .Z(n351) );
  XOR2_X1 U358 ( .A(KEYINPUT20), .B(n351), .Z(n309) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n307), .B(G120GAT), .ZN(n317) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(n317), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n533) );
  XOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .Z(n410) );
  XOR2_X1 U365 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n313) );
  NAND2_X1 U366 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XOR2_X1 U367 ( .A(n313), .B(n312), .Z(n316) );
  XOR2_X1 U368 ( .A(KEYINPUT71), .B(G64GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n396) );
  XNOR2_X1 U371 ( .A(n316), .B(n396), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n317), .B(KEYINPUT13), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(KEYINPUT33), .B(n320), .Z(n322) );
  XOR2_X1 U375 ( .A(G148GAT), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U376 ( .A(n439), .B(KEYINPUT70), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n410), .B(n323), .ZN(n324) );
  XNOR2_X1 U379 ( .A(G85GAT), .B(G92GAT), .ZN(n346) );
  XNOR2_X1 U380 ( .A(n324), .B(n346), .ZN(n579) );
  XNOR2_X1 U381 ( .A(KEYINPUT41), .B(n579), .ZN(n452) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n326) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U385 ( .A(n327), .B(KEYINPUT29), .Z(n335) );
  XOR2_X1 U386 ( .A(G113GAT), .B(G43GAT), .Z(n329) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(G29GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U389 ( .A(G8GAT), .B(KEYINPUT69), .Z(n331) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G197GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n341) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G50GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n348) );
  XOR2_X1 U397 ( .A(G1GAT), .B(KEYINPUT68), .Z(n339) );
  XNOR2_X1 U398 ( .A(G15GAT), .B(G22GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n375) );
  XOR2_X1 U400 ( .A(n348), .B(n375), .Z(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n576) );
  NAND2_X1 U402 ( .A1(n452), .A2(n576), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(KEYINPUT46), .ZN(n383) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n344) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(KEYINPUT66), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n350) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n345) );
  XOR2_X1 U408 ( .A(n350), .B(n349), .Z(n353) );
  XOR2_X1 U409 ( .A(G29GAT), .B(KEYINPUT74), .Z(n441) );
  XNOR2_X1 U410 ( .A(n351), .B(n441), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n361) );
  XOR2_X1 U412 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n355) );
  XNOR2_X1 U413 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT73), .B(G162GAT), .Z(n357) );
  XNOR2_X1 U416 ( .A(G190GAT), .B(G99GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n360) );
  XOR2_X1 U419 ( .A(G78GAT), .B(G211GAT), .Z(n363) );
  XNOR2_X1 U420 ( .A(G71GAT), .B(G155GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U422 ( .A(KEYINPUT79), .B(KEYINPUT13), .Z(n365) );
  XNOR2_X1 U423 ( .A(G57GAT), .B(G64GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U425 ( .A(n367), .B(n366), .Z(n372) );
  XOR2_X1 U426 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n369) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(KEYINPUT77), .B(n370), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n381) );
  XOR2_X1 U431 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n374) );
  XNOR2_X1 U432 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U434 ( .A(G8GAT), .B(KEYINPUT75), .Z(n395) );
  XOR2_X1 U435 ( .A(n395), .B(G127GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(n375), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(n379), .B(n378), .Z(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n491) );
  INV_X1 U440 ( .A(n491), .ZN(n583) );
  NOR2_X1 U441 ( .A1(n566), .A2(n583), .ZN(n382) );
  AND2_X1 U442 ( .A1(n383), .A2(n382), .ZN(n385) );
  INV_X1 U443 ( .A(KEYINPUT47), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n392) );
  INV_X1 U445 ( .A(KEYINPUT36), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n566), .B(n386), .ZN(n587) );
  NOR2_X1 U447 ( .A1(n491), .A2(n587), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n387), .B(KEYINPUT45), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n388), .A2(n579), .ZN(n389) );
  NOR2_X1 U450 ( .A1(n576), .A2(n389), .ZN(n390) );
  XNOR2_X1 U451 ( .A(KEYINPUT114), .B(n390), .ZN(n391) );
  NOR2_X1 U452 ( .A1(n392), .A2(n391), .ZN(n394) );
  XOR2_X1 U453 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n400) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G92GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U459 ( .A(n402), .B(n401), .Z(n408) );
  XNOR2_X1 U460 ( .A(n403), .B(KEYINPUT84), .ZN(n404) );
  XNOR2_X1 U461 ( .A(G197GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n296), .B(n405), .ZN(n417) );
  XNOR2_X1 U463 ( .A(n406), .B(n417), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n524) );
  NOR2_X1 U465 ( .A1(n532), .A2(n524), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n409), .B(KEYINPUT54), .ZN(n573) );
  XOR2_X1 U467 ( .A(n410), .B(KEYINPUT24), .Z(n412) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n413), .B(G204GAT), .Z(n416) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n415) );
  XNOR2_X1 U472 ( .A(G22GAT), .B(G148GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(n417), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT2), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U475 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U477 ( .A(G141GAT), .B(n422), .Z(n446) );
  XOR2_X1 U478 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n446), .B(n425), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n468) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G134GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(G120GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n435) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(KEYINPUT89), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n473) );
  INV_X1 U499 ( .A(n572), .ZN(n548) );
  NOR2_X1 U500 ( .A1(n468), .A2(n548), .ZN(n447) );
  AND2_X1 U501 ( .A1(n573), .A2(n447), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NOR2_X1 U503 ( .A1(n533), .A2(n449), .ZN(n451) );
  INV_X1 U504 ( .A(KEYINPUT119), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n565) );
  XNOR2_X1 U506 ( .A(n452), .B(KEYINPUT108), .ZN(n538) );
  NAND2_X1 U507 ( .A1(n565), .A2(n538), .ZN(n457) );
  XOR2_X1 U508 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n459) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT99), .B(n460), .Z(n481) );
  NAND2_X1 U515 ( .A1(n576), .A2(n579), .ZN(n494) );
  NOR2_X1 U516 ( .A1(n566), .A2(n491), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT16), .B(n461), .ZN(n479) );
  XNOR2_X1 U518 ( .A(KEYINPUT82), .B(n533), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n524), .B(KEYINPUT95), .ZN(n462) );
  XOR2_X1 U520 ( .A(n462), .B(KEYINPUT27), .Z(n471) );
  INV_X1 U521 ( .A(n528), .ZN(n515) );
  OR2_X1 U522 ( .A1(n471), .A2(n515), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n464), .A2(n535), .ZN(n476) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n467) );
  NOR2_X1 U525 ( .A1(n533), .A2(n524), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n468), .A2(n465), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n468), .A2(n533), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT96), .ZN(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT26), .B(n470), .ZN(n574) );
  OR2_X1 U531 ( .A1(n574), .A2(n471), .ZN(n547) );
  NAND2_X1 U532 ( .A1(n472), .A2(n547), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT98), .B(n477), .Z(n489) );
  INV_X1 U536 ( .A(n489), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n506) );
  NOR2_X1 U538 ( .A1(n494), .A2(n506), .ZN(n486) );
  NAND2_X1 U539 ( .A1(n486), .A2(n548), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  INV_X1 U541 ( .A(n524), .ZN(n510) );
  NAND2_X1 U542 ( .A1(n486), .A2(n510), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n484) );
  INV_X1 U545 ( .A(n533), .ZN(n512) );
  NAND2_X1 U546 ( .A1(n486), .A2(n512), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT103), .Z(n488) );
  NAND2_X1 U550 ( .A1(n486), .A2(n515), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n587), .A2(n489), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n491), .A2(n490), .ZN(n493) );
  NOR2_X1 U554 ( .A1(n522), .A2(n494), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n495), .Z(n504) );
  NOR2_X1 U556 ( .A1(n504), .A2(n572), .ZN(n499) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n524), .A2(n504), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n297), .ZN(G1329GAT) );
  XNOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n502) );
  NOR2_X1 U564 ( .A1(n533), .A2(n504), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n528), .A2(n504), .ZN(n505) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n508) );
  INV_X1 U570 ( .A(n576), .ZN(n550) );
  NAND2_X1 U571 ( .A1(n550), .A2(n538), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n521), .A2(n506), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n516), .A2(n548), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n510), .A2(n516), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n516), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(KEYINPUT110), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT111), .Z(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n572), .A2(n527), .ZN(n523) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n533), .A2(n527), .ZN(n526) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n550), .A2(n537), .ZN(n536) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  INV_X1 U602 ( .A(n537), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n543), .A2(n538), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n543), .A2(n583), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U609 ( .A1(n543), .A2(n566), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n532), .A2(n547), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n552) );
  NOR2_X1 U614 ( .A1(n550), .A2(n552), .ZN(n551) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n554) );
  INV_X1 U617 ( .A(n552), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n559), .A2(n452), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(n555), .B(KEYINPUT52), .Z(n557) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n583), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n576), .A2(n565), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n583), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(n571), .Z(n578) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n584), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n581) );
  INV_X1 U645 ( .A(n584), .ZN(n586) );
  OR2_X1 U646 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

