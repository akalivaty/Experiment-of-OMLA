

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758;

  OR2_X1 U375 ( .A1(n562), .A2(n563), .ZN(n651) );
  NAND2_X1 U376 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U377 ( .A(n367), .B(n484), .ZN(n725) );
  XNOR2_X1 U378 ( .A(n380), .B(G146), .ZN(n518) );
  XNOR2_X1 U379 ( .A(n741), .B(G101), .ZN(n380) );
  XNOR2_X1 U380 ( .A(n515), .B(n468), .ZN(n738) );
  BUF_X1 U381 ( .A(G128), .Z(n352) );
  INV_X2 U382 ( .A(G128), .ZN(n425) );
  AND2_X2 U383 ( .A1(n460), .A2(n364), .ZN(n417) );
  AND2_X1 U384 ( .A1(n662), .A2(n386), .ZN(n615) );
  INV_X2 U385 ( .A(G953), .ZN(n749) );
  XNOR2_X2 U386 ( .A(n455), .B(G107), .ZN(n544) );
  XNOR2_X2 U387 ( .A(G116), .B(G122), .ZN(n455) );
  NOR2_X2 U388 ( .A1(n619), .A2(n620), .ZN(n418) );
  XNOR2_X2 U389 ( .A(n496), .B(n385), .ZN(n384) );
  XNOR2_X2 U390 ( .A(n421), .B(n434), .ZN(n662) );
  XNOR2_X2 U391 ( .A(n591), .B(n355), .ZN(n676) );
  NAND2_X1 U392 ( .A1(n431), .A2(n444), .ZN(n403) );
  XNOR2_X1 U393 ( .A(n404), .B(n446), .ZN(n431) );
  NOR2_X2 U394 ( .A1(n435), .A2(n753), .ZN(n622) );
  XNOR2_X1 U395 ( .A(n569), .B(KEYINPUT32), .ZN(n458) );
  NAND2_X1 U396 ( .A1(n374), .A2(n371), .ZN(n653) );
  XNOR2_X1 U397 ( .A(n612), .B(n611), .ZN(n755) );
  NAND2_X1 U398 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U399 ( .A(n394), .B(n361), .ZN(n609) );
  XNOR2_X1 U400 ( .A(n489), .B(KEYINPUT19), .ZN(n587) );
  BUF_X1 U401 ( .A(n575), .Z(n421) );
  INV_X1 U402 ( .A(KEYINPUT107), .ZN(n611) );
  AND2_X1 U403 ( .A1(n629), .A2(n628), .ZN(n720) );
  XNOR2_X1 U404 ( .A(n415), .B(n518), .ZN(n710) );
  AND2_X1 U405 ( .A1(n457), .A2(n458), .ZN(n573) );
  XNOR2_X1 U406 ( .A(G902), .B(KEYINPUT15), .ZN(n624) );
  XOR2_X1 U407 ( .A(G137), .B(G140), .Z(n494) );
  XNOR2_X1 U408 ( .A(n433), .B(G104), .ZN(n533) );
  INV_X1 U409 ( .A(G113), .ZN(n433) );
  XNOR2_X1 U410 ( .A(n426), .B(G472), .ZN(n556) );
  OR2_X1 U411 ( .A1(n635), .A2(G902), .ZN(n426) );
  NAND2_X1 U412 ( .A1(n587), .A2(n490), .ZN(n464) );
  INV_X1 U413 ( .A(KEYINPUT0), .ZN(n463) );
  XNOR2_X1 U414 ( .A(n382), .B(n381), .ZN(n505) );
  NOR2_X1 U415 ( .A1(n722), .A2(G902), .ZN(n506) );
  XNOR2_X1 U416 ( .A(n504), .B(KEYINPUT91), .ZN(n381) );
  INV_X1 U417 ( .A(G134), .ZN(n469) );
  AND2_X1 U418 ( .A1(n636), .A2(n564), .ZN(n571) );
  NAND2_X1 U419 ( .A1(n653), .A2(n639), .ZN(n378) );
  NOR2_X1 U420 ( .A1(n580), .A2(n691), .ZN(n596) );
  OR2_X1 U421 ( .A1(G237), .A2(G902), .ZN(n488) );
  INV_X1 U422 ( .A(KEYINPUT10), .ZN(n385) );
  XNOR2_X1 U423 ( .A(G140), .B(KEYINPUT93), .ZN(n526) );
  NAND2_X1 U424 ( .A1(n624), .A2(KEYINPUT79), .ZN(n461) );
  INV_X1 U425 ( .A(n494), .ZN(n468) );
  XNOR2_X1 U426 ( .A(G104), .B(G107), .ZN(n493) );
  XOR2_X1 U427 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n479) );
  XOR2_X1 U428 ( .A(KEYINPUT69), .B(G110), .Z(n491) );
  NOR2_X1 U429 ( .A1(n445), .A2(n659), .ZN(n444) );
  INV_X1 U430 ( .A(n657), .ZN(n445) );
  INV_X1 U431 ( .A(n576), .ZN(n396) );
  XNOR2_X1 U432 ( .A(KEYINPUT38), .B(KEYINPUT71), .ZN(n434) );
  NAND2_X1 U433 ( .A1(n588), .A2(n430), .ZN(n429) );
  INV_X1 U434 ( .A(n589), .ZN(n430) );
  XNOR2_X1 U435 ( .A(n540), .B(n539), .ZN(n560) );
  XNOR2_X1 U436 ( .A(n556), .B(KEYINPUT6), .ZN(n576) );
  XNOR2_X1 U437 ( .A(n544), .B(n456), .ZN(n367) );
  INV_X1 U438 ( .A(n533), .ZN(n456) );
  XNOR2_X1 U439 ( .A(n523), .B(n522), .ZN(n467) );
  XNOR2_X1 U440 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X1 U441 ( .A(n511), .B(n471), .ZN(n517) );
  NAND2_X1 U442 ( .A1(n365), .A2(G472), .ZN(n454) );
  NAND2_X1 U443 ( .A1(n359), .A2(n676), .ZN(n457) );
  INV_X1 U444 ( .A(KEYINPUT70), .ZN(n406) );
  INV_X1 U445 ( .A(KEYINPUT68), .ZN(n423) );
  INV_X1 U446 ( .A(KEYINPUT104), .ZN(n443) );
  NAND2_X1 U447 ( .A1(G953), .A2(G902), .ZN(n577) );
  XOR2_X1 U448 ( .A(KEYINPUT96), .B(KEYINPUT94), .Z(n530) );
  XOR2_X1 U449 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n527) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n446) );
  NOR2_X1 U451 ( .A1(n675), .A2(n443), .ZN(n438) );
  XNOR2_X1 U452 ( .A(n503), .B(n502), .ZN(n507) );
  XNOR2_X1 U453 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n502) );
  XOR2_X1 U454 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n504) );
  NAND2_X1 U455 ( .A1(n507), .A2(G217), .ZN(n382) );
  INV_X1 U456 ( .A(KEYINPUT67), .ZN(n470) );
  NOR2_X1 U457 ( .A1(G953), .A2(G237), .ZN(n528) );
  NAND2_X1 U458 ( .A1(n571), .A2(n409), .ZN(n572) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n409) );
  INV_X1 U460 ( .A(KEYINPUT83), .ZN(n400) );
  XOR2_X1 U461 ( .A(KEYINPUT3), .B(G119), .Z(n509) );
  NAND2_X1 U462 ( .A1(n662), .A2(n661), .ZN(n387) );
  NOR2_X1 U463 ( .A1(n676), .A2(n675), .ZN(n557) );
  XNOR2_X1 U464 ( .A(G137), .B(KEYINPUT72), .ZN(n512) );
  XOR2_X1 U465 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n513) );
  XNOR2_X1 U466 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U467 ( .A(G113), .B(G116), .ZN(n510) );
  XNOR2_X1 U468 ( .A(n384), .B(n356), .ZN(n499) );
  XNOR2_X1 U469 ( .A(n352), .B(G110), .ZN(n495) );
  XOR2_X1 U470 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n542) );
  XNOR2_X1 U471 ( .A(G134), .B(KEYINPUT9), .ZN(n541) );
  XNOR2_X1 U472 ( .A(n414), .B(n383), .ZN(n397) );
  AND2_X1 U473 ( .A1(n733), .A2(n353), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n407), .B(n419), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n492), .B(n493), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n366), .B(n485), .ZN(n705) );
  XNOR2_X1 U477 ( .A(n725), .B(n491), .ZN(n366) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n475) );
  XNOR2_X1 U479 ( .A(n520), .B(KEYINPUT33), .ZN(n670) );
  NAND2_X1 U480 ( .A1(n557), .A2(n396), .ZN(n520) );
  NOR2_X1 U481 ( .A1(n651), .A2(n395), .ZN(n608) );
  NAND2_X1 U482 ( .A1(n396), .A2(n583), .ZN(n395) );
  XNOR2_X1 U483 ( .A(n615), .B(n614), .ZN(n686) );
  NOR2_X1 U484 ( .A1(n664), .A2(n581), .ZN(n386) );
  NAND2_X1 U485 ( .A1(n608), .A2(n421), .ZN(n394) );
  NAND2_X1 U486 ( .A1(n684), .A2(n377), .ZN(n375) );
  INV_X1 U487 ( .A(n558), .ZN(n373) );
  INV_X1 U488 ( .A(KEYINPUT28), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n555), .B(n402), .ZN(n401) );
  INV_X1 U490 ( .A(KEYINPUT22), .ZN(n402) );
  INV_X1 U491 ( .A(n565), .ZN(n679) );
  AND2_X1 U492 ( .A1(n401), .A2(n576), .ZN(n568) );
  XNOR2_X1 U493 ( .A(n450), .B(n447), .ZN(n722) );
  XNOR2_X1 U494 ( .A(n449), .B(n448), .ZN(n447) );
  XNOR2_X1 U495 ( .A(n499), .B(n500), .ZN(n450) );
  XNOR2_X1 U496 ( .A(n498), .B(n354), .ZN(n448) );
  XNOR2_X1 U497 ( .A(n552), .B(KEYINPUT35), .ZN(n465) );
  NAND2_X1 U498 ( .A1(n467), .A2(n604), .ZN(n466) );
  INV_X1 U499 ( .A(KEYINPUT82), .ZN(n552) );
  NAND2_X1 U500 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U501 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X1 U502 ( .A1(n684), .A2(n377), .ZN(n372) );
  NAND2_X1 U503 ( .A1(n568), .A2(n408), .ZN(n636) );
  AND2_X1 U504 ( .A1(n676), .A2(n410), .ZN(n408) );
  XNOR2_X1 U505 ( .A(n454), .B(n363), .ZN(n453) );
  INV_X1 U506 ( .A(KEYINPUT60), .ZN(n411) );
  INV_X1 U507 ( .A(n457), .ZN(n643) );
  INV_X1 U508 ( .A(n676), .ZN(n610) );
  AND2_X1 U509 ( .A1(n501), .A2(n462), .ZN(n353) );
  XOR2_X1 U510 ( .A(G119), .B(KEYINPUT88), .Z(n354) );
  XOR2_X1 U511 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n355) );
  XOR2_X1 U512 ( .A(KEYINPUT78), .B(KEYINPUT89), .Z(n356) );
  OR2_X1 U513 ( .A1(n574), .A2(KEYINPUT44), .ZN(n357) );
  AND2_X1 U514 ( .A1(n439), .A2(n436), .ZN(n358) );
  AND2_X1 U515 ( .A1(n566), .A2(n565), .ZN(n359) );
  AND2_X1 U516 ( .A1(n405), .A2(n595), .ZN(n360) );
  XOR2_X1 U517 ( .A(KEYINPUT36), .B(KEYINPUT84), .Z(n361) );
  XOR2_X1 U518 ( .A(n463), .B(KEYINPUT85), .Z(n362) );
  XOR2_X1 U519 ( .A(n635), .B(KEYINPUT62), .Z(n363) );
  INV_X1 U520 ( .A(n624), .ZN(n501) );
  AND2_X1 U521 ( .A1(n626), .A2(n461), .ZN(n364) );
  NOR2_X1 U522 ( .A1(G952), .A2(n749), .ZN(n724) );
  INV_X1 U523 ( .A(n724), .ZN(n452) );
  AND2_X2 U524 ( .A1(n629), .A2(n628), .ZN(n365) );
  NAND2_X1 U525 ( .A1(n417), .A2(n459), .ZN(n629) );
  INV_X1 U526 ( .A(n591), .ZN(n439) );
  NAND2_X1 U527 ( .A1(n368), .A2(n572), .ZN(n370) );
  NAND2_X1 U528 ( .A1(n570), .A2(n573), .ZN(n368) );
  NAND2_X1 U529 ( .A1(n369), .A2(n357), .ZN(n399) );
  XNOR2_X1 U530 ( .A(n370), .B(n400), .ZN(n369) );
  NAND2_X1 U531 ( .A1(n558), .A2(n377), .ZN(n376) );
  INV_X1 U532 ( .A(KEYINPUT31), .ZN(n377) );
  NAND2_X1 U533 ( .A1(n378), .A2(n592), .ZN(n564) );
  XNOR2_X2 U534 ( .A(n379), .B(G469), .ZN(n591) );
  NOR2_X2 U535 ( .A1(n710), .A2(G902), .ZN(n379) );
  XNOR2_X1 U536 ( .A(n380), .B(n483), .ZN(n485) );
  INV_X1 U537 ( .A(n384), .ZN(n383) );
  XNOR2_X1 U538 ( .A(n384), .B(n738), .ZN(n739) );
  NOR2_X1 U539 ( .A1(n665), .A2(n387), .ZN(n666) );
  NAND2_X1 U540 ( .A1(n388), .A2(n423), .ZN(n392) );
  NAND2_X1 U541 ( .A1(n389), .A2(n360), .ZN(n388) );
  INV_X1 U542 ( .A(n393), .ZN(n389) );
  NAND2_X1 U543 ( .A1(n613), .A2(n755), .ZN(n393) );
  NAND2_X1 U544 ( .A1(n392), .A2(n390), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n391), .A2(n360), .ZN(n390) );
  NOR2_X1 U546 ( .A1(n393), .A2(n423), .ZN(n391) );
  NOR2_X1 U547 ( .A1(n630), .A2(G902), .ZN(n540) );
  XNOR2_X1 U548 ( .A(n398), .B(n397), .ZN(n630) );
  XNOR2_X1 U549 ( .A(n534), .B(n535), .ZN(n398) );
  XNOR2_X2 U550 ( .A(n399), .B(KEYINPUT45), .ZN(n733) );
  AND2_X1 U551 ( .A1(n401), .A2(n588), .ZN(n566) );
  XNOR2_X2 U552 ( .A(n403), .B(KEYINPUT81), .ZN(n748) );
  NOR2_X1 U553 ( .A1(n627), .A2(n403), .ZN(n700) );
  NAND2_X1 U554 ( .A1(n432), .A2(n422), .ZN(n404) );
  XNOR2_X1 U555 ( .A(n594), .B(n406), .ZN(n405) );
  XNOR2_X1 U556 ( .A(n428), .B(n427), .ZN(n590) );
  AND2_X1 U557 ( .A1(n442), .A2(n441), .ZN(n440) );
  INV_X1 U558 ( .A(n738), .ZN(n407) );
  XNOR2_X1 U559 ( .A(n518), .B(n519), .ZN(n635) );
  BUF_X1 U560 ( .A(n673), .Z(n410) );
  NAND2_X1 U561 ( .A1(n591), .A2(n443), .ZN(n442) );
  NOR2_X1 U562 ( .A1(n619), .A2(n602), .ZN(n603) );
  NAND2_X1 U563 ( .A1(n575), .A2(n661), .ZN(n489) );
  XNOR2_X1 U564 ( .A(n487), .B(n486), .ZN(n575) );
  NAND2_X1 U565 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U566 ( .A(n621), .B(KEYINPUT40), .ZN(n435) );
  NAND2_X1 U567 ( .A1(n675), .A2(n443), .ZN(n441) );
  XNOR2_X1 U568 ( .A(n412), .B(n411), .ZN(G60) );
  NAND2_X1 U569 ( .A1(n416), .A2(n452), .ZN(n412) );
  XNOR2_X1 U570 ( .A(n418), .B(KEYINPUT39), .ZN(n623) );
  NAND2_X1 U571 ( .A1(n546), .A2(G221), .ZN(n449) );
  INV_X1 U572 ( .A(n521), .ZN(n558) );
  NAND2_X1 U573 ( .A1(n521), .A2(n554), .ZN(n555) );
  XNOR2_X2 U574 ( .A(n464), .B(n362), .ZN(n521) );
  XNOR2_X1 U575 ( .A(n413), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U576 ( .A1(n709), .A2(n724), .ZN(n413) );
  XNOR2_X1 U577 ( .A(n533), .B(KEYINPUT95), .ZN(n414) );
  XNOR2_X2 U578 ( .A(n506), .B(n505), .ZN(n673) );
  XNOR2_X1 U579 ( .A(n634), .B(n633), .ZN(n416) );
  NAND2_X1 U580 ( .A1(n365), .A2(G475), .ZN(n634) );
  NAND2_X1 U581 ( .A1(n420), .A2(n748), .ZN(n459) );
  NAND2_X1 U582 ( .A1(n733), .A2(KEYINPUT2), .ZN(n627) );
  XNOR2_X2 U583 ( .A(n545), .B(n424), .ZN(n741) );
  INV_X1 U584 ( .A(n477), .ZN(n424) );
  XNOR2_X2 U585 ( .A(n425), .B(G143), .ZN(n545) );
  NOR2_X1 U586 ( .A1(n565), .A2(n429), .ZN(n428) );
  XNOR2_X1 U587 ( .A(n622), .B(KEYINPUT46), .ZN(n432) );
  XNOR2_X1 U588 ( .A(n435), .B(n754), .ZN(G33) );
  INV_X1 U589 ( .A(n675), .ZN(n436) );
  NAND2_X1 U590 ( .A1(n440), .A2(n437), .ZN(n597) );
  NAND2_X1 U591 ( .A1(n439), .A2(n438), .ZN(n437) );
  XNOR2_X1 U592 ( .A(n451), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U593 ( .A(G146), .B(G125), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n458), .B(G119), .ZN(G21) );
  NAND2_X1 U595 ( .A1(n733), .A2(n748), .ZN(n698) );
  NAND2_X1 U596 ( .A1(n698), .A2(KEYINPUT79), .ZN(n460) );
  INV_X1 U597 ( .A(KEYINPUT79), .ZN(n462) );
  XNOR2_X2 U598 ( .A(n466), .B(n465), .ZN(n758) );
  XNOR2_X2 U599 ( .A(n524), .B(n469), .ZN(n515) );
  XNOR2_X2 U600 ( .A(n470), .B(G131), .ZN(n524) );
  AND2_X1 U601 ( .A1(n528), .A2(G210), .ZN(n471) );
  AND2_X1 U602 ( .A1(G227), .A2(n749), .ZN(n472) );
  XOR2_X1 U603 ( .A(n707), .B(n706), .Z(n473) );
  INV_X1 U604 ( .A(KEYINPUT76), .ZN(n606) );
  XNOR2_X1 U605 ( .A(n496), .B(n480), .ZN(n481) );
  XNOR2_X1 U606 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U607 ( .A(n491), .B(n472), .ZN(n492) );
  INV_X1 U608 ( .A(n672), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n515), .B(n514), .ZN(n516) );
  AND2_X1 U610 ( .A1(n588), .A2(n582), .ZN(n583) );
  NOR2_X1 U611 ( .A1(n664), .A2(n553), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n517), .B(n516), .ZN(n519) );
  INV_X1 U613 ( .A(n700), .ZN(n628) );
  XNOR2_X1 U614 ( .A(n598), .B(KEYINPUT73), .ZN(n601) );
  AND2_X1 U615 ( .A1(n610), .A2(n588), .ZN(n567) );
  XNOR2_X1 U616 ( .A(n708), .B(n473), .ZN(n709) );
  OR2_X1 U617 ( .A1(n623), .A2(n654), .ZN(n657) );
  INV_X1 U618 ( .A(G952), .ZN(n692) );
  NOR2_X1 U619 ( .A1(G953), .A2(n692), .ZN(n579) );
  NOR2_X1 U620 ( .A1(G898), .A2(n577), .ZN(n474) );
  NOR2_X1 U621 ( .A1(n579), .A2(n474), .ZN(n476) );
  XOR2_X1 U622 ( .A(KEYINPUT14), .B(n475), .Z(n691) );
  NOR2_X1 U623 ( .A1(n476), .A2(n691), .ZN(n490) );
  XNOR2_X1 U624 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n477) );
  NAND2_X1 U625 ( .A1(G224), .A2(n749), .ZN(n478) );
  XNOR2_X1 U626 ( .A(n479), .B(n478), .ZN(n482) );
  XOR2_X1 U627 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n480) );
  XNOR2_X1 U628 ( .A(n509), .B(KEYINPUT16), .ZN(n484) );
  NOR2_X1 U629 ( .A1(n705), .A2(n501), .ZN(n487) );
  NAND2_X1 U630 ( .A1(G210), .A2(n488), .ZN(n486) );
  NAND2_X1 U631 ( .A1(n488), .A2(G214), .ZN(n661) );
  XNOR2_X1 U632 ( .A(n495), .B(n494), .ZN(n500) );
  NAND2_X1 U633 ( .A1(G234), .A2(n749), .ZN(n497) );
  XOR2_X1 U634 ( .A(KEYINPUT8), .B(n497), .Z(n546) );
  XOR2_X1 U635 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n498) );
  NAND2_X1 U636 ( .A1(n624), .A2(G234), .ZN(n503) );
  NAND2_X1 U637 ( .A1(n507), .A2(G221), .ZN(n508) );
  XOR2_X1 U638 ( .A(KEYINPUT21), .B(n508), .Z(n672) );
  XNOR2_X1 U639 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U640 ( .A1(n521), .A2(n670), .ZN(n523) );
  XNOR2_X1 U641 ( .A(n524), .B(G143), .ZN(n525) );
  XNOR2_X1 U642 ( .A(n525), .B(G122), .ZN(n535) );
  XNOR2_X1 U643 ( .A(n527), .B(n526), .ZN(n532) );
  NAND2_X1 U644 ( .A1(G214), .A2(n528), .ZN(n529) );
  XNOR2_X1 U645 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U646 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U647 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n537) );
  XNOR2_X1 U648 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n536) );
  XNOR2_X1 U649 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U650 ( .A(G475), .B(n538), .ZN(n539) );
  XNOR2_X1 U651 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n544), .B(n543), .ZN(n550) );
  XOR2_X1 U653 ( .A(n545), .B(KEYINPUT101), .Z(n548) );
  NAND2_X1 U654 ( .A1(G217), .A2(n546), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U656 ( .A(n550), .B(n549), .ZN(n716) );
  NOR2_X1 U657 ( .A1(n716), .A2(G902), .ZN(n551) );
  XNOR2_X1 U658 ( .A(n551), .B(G478), .ZN(n561) );
  NOR2_X1 U659 ( .A1(n560), .A2(n561), .ZN(n604) );
  NAND2_X1 U660 ( .A1(n560), .A2(n561), .ZN(n664) );
  INV_X1 U661 ( .A(n556), .ZN(n565) );
  NAND2_X1 U662 ( .A1(n679), .A2(n557), .ZN(n684) );
  NOR2_X1 U663 ( .A1(n679), .A2(n558), .ZN(n559) );
  NAND2_X1 U664 ( .A1(n358), .A2(n559), .ZN(n639) );
  XNOR2_X1 U665 ( .A(n560), .B(KEYINPUT100), .ZN(n562) );
  INV_X1 U666 ( .A(n561), .ZN(n563) );
  NAND2_X1 U667 ( .A1(n563), .A2(n562), .ZN(n654) );
  NAND2_X1 U668 ( .A1(n651), .A2(n654), .ZN(n592) );
  AND2_X1 U669 ( .A1(n571), .A2(n758), .ZN(n570) );
  INV_X1 U670 ( .A(n673), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U672 ( .A1(n758), .A2(n573), .ZN(n574) );
  XOR2_X1 U673 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n585) );
  INV_X1 U674 ( .A(n661), .ZN(n581) );
  NOR2_X1 U675 ( .A1(G900), .A2(n577), .ZN(n578) );
  NOR2_X1 U676 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U677 ( .A1(n596), .A2(n672), .ZN(n589) );
  NOR2_X1 U678 ( .A1(n581), .A2(n589), .ZN(n582) );
  NAND2_X1 U679 ( .A1(n608), .A2(n676), .ZN(n584) );
  XOR2_X1 U680 ( .A(n585), .B(n584), .Z(n586) );
  NOR2_X1 U681 ( .A1(n421), .A2(n586), .ZN(n659) );
  NOR2_X1 U682 ( .A1(n591), .A2(n590), .ZN(n616) );
  NAND2_X1 U683 ( .A1(n587), .A2(n616), .ZN(n648) );
  INV_X1 U684 ( .A(n592), .ZN(n665) );
  OR2_X1 U685 ( .A1(KEYINPUT47), .A2(n665), .ZN(n593) );
  NOR2_X1 U686 ( .A1(n648), .A2(n593), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n648), .A2(KEYINPUT47), .ZN(n595) );
  INV_X1 U688 ( .A(n421), .ZN(n602) );
  NAND2_X1 U689 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U690 ( .A1(n556), .A2(n661), .ZN(n599) );
  XOR2_X1 U691 ( .A(KEYINPUT30), .B(n599), .Z(n600) );
  NAND2_X1 U692 ( .A1(n601), .A2(n600), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n604), .A2(n603), .ZN(n647) );
  NAND2_X1 U694 ( .A1(KEYINPUT47), .A2(n665), .ZN(n605) );
  NAND2_X1 U695 ( .A1(n647), .A2(n605), .ZN(n607) );
  XNOR2_X1 U696 ( .A(n607), .B(n606), .ZN(n613) );
  XOR2_X1 U697 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n618) );
  XNOR2_X1 U698 ( .A(KEYINPUT41), .B(KEYINPUT105), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n686), .A2(n616), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n618), .B(n617), .ZN(n753) );
  INV_X1 U701 ( .A(n662), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n623), .A2(n651), .ZN(n621) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n697) );
  XNOR2_X1 U704 ( .A(KEYINPUT80), .B(n624), .ZN(n625) );
  OR2_X1 U705 ( .A1(n697), .A2(n625), .ZN(n626) );
  XNOR2_X1 U706 ( .A(KEYINPUT118), .B(KEYINPUT59), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT66), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U709 ( .A(n636), .ZN(n637) );
  XOR2_X1 U710 ( .A(G101), .B(n637), .Z(G3) );
  NOR2_X1 U711 ( .A1(n651), .A2(n639), .ZN(n638) );
  XOR2_X1 U712 ( .A(G104), .B(n638), .Z(G6) );
  NOR2_X1 U713 ( .A1(n654), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U716 ( .A(G107), .B(n642), .ZN(G9) );
  XOR2_X1 U717 ( .A(G110), .B(n643), .Z(G12) );
  NOR2_X1 U718 ( .A1(n654), .A2(n648), .ZN(n645) );
  XNOR2_X1 U719 ( .A(KEYINPUT29), .B(KEYINPUT108), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n352), .B(n646), .ZN(G30) );
  XNOR2_X1 U722 ( .A(G143), .B(n647), .ZN(G45) );
  NOR2_X1 U723 ( .A1(n651), .A2(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(G146), .B(KEYINPUT109), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(G48) );
  NOR2_X1 U726 ( .A1(n651), .A2(n653), .ZN(n652) );
  XOR2_X1 U727 ( .A(G113), .B(n652), .Z(G15) );
  NOR2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT110), .B(n655), .Z(n656) );
  XNOR2_X1 U730 ( .A(G116), .B(n656), .ZN(G18) );
  XNOR2_X1 U731 ( .A(G134), .B(KEYINPUT112), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(G36) );
  XNOR2_X1 U733 ( .A(G140), .B(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(KEYINPUT113), .ZN(G42) );
  NAND2_X1 U735 ( .A1(n686), .A2(n670), .ZN(n696) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(n666), .Z(n667) );
  NOR2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U740 ( .A(KEYINPUT116), .B(n669), .Z(n671) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n689) );
  NOR2_X1 U742 ( .A1(n410), .A2(n672), .ZN(n674) );
  XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n674), .ZN(n682) );
  XOR2_X1 U744 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n678) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT51), .B(n685), .Z(n687) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U753 ( .A(KEYINPUT52), .B(n690), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n702) );
  AND2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n749), .A2(n703), .ZN(n704) );
  XOR2_X1 U761 ( .A(KEYINPUT53), .B(n704), .Z(G75) );
  NAND2_X1 U762 ( .A1(n720), .A2(G210), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT77), .B(KEYINPUT55), .Z(n707) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT54), .ZN(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n710), .B(KEYINPUT57), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U768 ( .A1(n365), .A2(G469), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n724), .A2(n715), .ZN(G54) );
  XOR2_X1 U771 ( .A(n716), .B(KEYINPUT119), .Z(n718) );
  NAND2_X1 U772 ( .A1(n365), .A2(G478), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n724), .A2(n719), .ZN(G63) );
  NAND2_X1 U775 ( .A1(G217), .A2(n365), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(G66) );
  XNOR2_X1 U778 ( .A(n725), .B(G110), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n726), .B(KEYINPUT121), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n727), .B(G101), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n749), .A2(G898), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n737) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n731), .A2(G898), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n732), .B(KEYINPUT120), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n733), .A2(n749), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(G69) );
  XNOR2_X1 U790 ( .A(KEYINPUT122), .B(n739), .ZN(n740) );
  XOR2_X1 U791 ( .A(n741), .B(n740), .Z(n747) );
  XOR2_X1 U792 ( .A(n747), .B(G227), .Z(n742) );
  XNOR2_X1 U793 ( .A(n742), .B(KEYINPUT123), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n743), .A2(G900), .ZN(n744) );
  XOR2_X1 U795 ( .A(KEYINPUT124), .B(n744), .Z(n745) );
  NOR2_X1 U796 ( .A1(n749), .A2(n745), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(KEYINPUT125), .ZN(n752) );
  XOR2_X1 U798 ( .A(n748), .B(n747), .Z(n750) );
  NAND2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U801 ( .A(n753), .B(G137), .Z(G39) );
  XOR2_X1 U802 ( .A(G131), .B(KEYINPUT126), .Z(n754) );
  XNOR2_X1 U803 ( .A(KEYINPUT37), .B(KEYINPUT111), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U805 ( .A(G125), .B(n757), .ZN(G27) );
  XNOR2_X1 U806 ( .A(G122), .B(n758), .ZN(G24) );
endmodule

