

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U326 ( .A(n328), .B(n327), .Z(n293) );
  NOR2_X1 U327 ( .A1(n510), .A2(n508), .ZN(n466) );
  XNOR2_X1 U328 ( .A(n295), .B(KEYINPUT80), .ZN(n296) );
  XNOR2_X1 U329 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U330 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U331 ( .A(n329), .B(n293), .ZN(n330) );
  XNOR2_X1 U332 ( .A(n312), .B(n311), .ZN(n584) );
  OR2_X1 U333 ( .A1(n532), .A2(n496), .ZN(n485) );
  NOR2_X1 U334 ( .A1(n510), .A2(n461), .ZN(n574) );
  XNOR2_X1 U335 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U336 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  XNOR2_X1 U338 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  XNOR2_X1 U339 ( .A(G71GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n294), .B(KEYINPUT13), .ZN(n370) );
  XOR2_X1 U341 ( .A(G106GAT), .B(G78GAT), .Z(n451) );
  XOR2_X1 U342 ( .A(n370), .B(n451), .Z(n297) );
  NAND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G148GAT), .Z(n422) );
  XOR2_X1 U345 ( .A(n422), .B(KEYINPUT33), .Z(n299) );
  NAND2_X1 U346 ( .A1(n298), .A2(n299), .ZN(n303) );
  INV_X1 U347 ( .A(n298), .ZN(n301) );
  INV_X1 U348 ( .A(n299), .ZN(n300) );
  NAND2_X1 U349 ( .A1(n301), .A2(n300), .ZN(n302) );
  NAND2_X1 U350 ( .A1(n303), .A2(n302), .ZN(n312) );
  XOR2_X1 U351 ( .A(G64GAT), .B(G92GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(G176GAT), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n339) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .ZN(n306) );
  XOR2_X1 U355 ( .A(n306), .B(KEYINPUT79), .Z(n407) );
  XOR2_X1 U356 ( .A(n339), .B(n407), .Z(n310) );
  XOR2_X1 U357 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n308) );
  XNOR2_X1 U358 ( .A(KEYINPUT78), .B(KEYINPUT31), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  INV_X1 U360 ( .A(KEYINPUT41), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n584), .B(n313), .ZN(n367) );
  XNOR2_X1 U362 ( .A(KEYINPUT112), .B(n367), .ZN(n548) );
  XOR2_X1 U363 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n315) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n333) );
  INV_X1 U366 ( .A(KEYINPUT17), .ZN(n316) );
  NAND2_X1 U367 ( .A1(KEYINPUT19), .A2(n316), .ZN(n319) );
  INV_X1 U368 ( .A(KEYINPUT19), .ZN(n317) );
  NAND2_X1 U369 ( .A1(n317), .A2(KEYINPUT17), .ZN(n318) );
  NAND2_X1 U370 ( .A1(n319), .A2(n318), .ZN(n321) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n344) );
  XOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT0), .Z(n427) );
  XNOR2_X1 U374 ( .A(n344), .B(n427), .ZN(n323) );
  XOR2_X1 U375 ( .A(G43GAT), .B(G190GAT), .Z(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G71GAT), .Z(n325) );
  XNOR2_X1 U378 ( .A(G15GAT), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(n326), .ZN(n329) );
  XOR2_X1 U381 ( .A(G127GAT), .B(G120GAT), .Z(n328) );
  NAND2_X1 U382 ( .A1(G227GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U383 ( .A(n333), .B(n332), .Z(n545) );
  INV_X1 U384 ( .A(n545), .ZN(n510) );
  XOR2_X1 U385 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n335) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U388 ( .A(n336), .B(KEYINPUT99), .Z(n338) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XOR2_X1 U390 ( .A(G8GAT), .B(G183GAT), .Z(n373) );
  XNOR2_X1 U391 ( .A(n398), .B(n373), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U394 ( .A(KEYINPUT91), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U395 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(G197GAT), .B(n343), .Z(n459) );
  XNOR2_X1 U398 ( .A(n344), .B(n459), .ZN(n345) );
  XOR2_X1 U399 ( .A(n346), .B(n345), .Z(n536) );
  INV_X1 U400 ( .A(n536), .ZN(n508) );
  XOR2_X1 U401 ( .A(KEYINPUT120), .B(KEYINPUT46), .Z(n369) );
  XOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n348) );
  XNOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U405 ( .A(G8GAT), .B(G197GAT), .Z(n350) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U409 ( .A(G50GAT), .B(G141GAT), .Z(n442) );
  XNOR2_X1 U410 ( .A(G29GAT), .B(G113GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n353), .B(G1GAT), .ZN(n426) );
  XOR2_X1 U412 ( .A(n442), .B(n426), .Z(n355) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT69), .B(KEYINPUT75), .Z(n357) );
  XNOR2_X1 U416 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U419 ( .A(G43GAT), .B(KEYINPUT7), .Z(n361) );
  XNOR2_X1 U420 ( .A(KEYINPUT73), .B(KEYINPUT8), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n406) );
  XNOR2_X1 U422 ( .A(G15GAT), .B(G22GAT), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n362), .B(KEYINPUT74), .ZN(n375) );
  XNOR2_X1 U424 ( .A(n406), .B(n375), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U426 ( .A(n366), .B(n365), .Z(n518) );
  INV_X1 U427 ( .A(n518), .ZN(n580) );
  NAND2_X1 U428 ( .A1(n580), .A2(n367), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n386) );
  XOR2_X1 U430 ( .A(n370), .B(KEYINPUT12), .Z(n372) );
  NAND2_X1 U431 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U433 ( .A(n374), .B(n373), .Z(n377) );
  XOR2_X1 U434 ( .A(G127GAT), .B(G155GAT), .Z(n421) );
  XNOR2_X1 U435 ( .A(n375), .B(n421), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G78GAT), .Z(n379) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT86), .Z(n381) );
  XNOR2_X1 U441 ( .A(KEYINPUT85), .B(KEYINPUT14), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U443 ( .A(n383), .B(n382), .Z(n384) );
  XOR2_X1 U444 ( .A(n385), .B(n384), .Z(n588) );
  XOR2_X1 U445 ( .A(KEYINPUT119), .B(n588), .Z(n571) );
  NOR2_X1 U446 ( .A1(n386), .A2(n571), .ZN(n409) );
  XOR2_X1 U447 ( .A(KEYINPUT83), .B(KEYINPUT65), .Z(n388) );
  XNOR2_X1 U448 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U450 ( .A(KEYINPUT82), .B(KEYINPUT67), .Z(n390) );
  XNOR2_X1 U451 ( .A(G50GAT), .B(G92GAT), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U453 ( .A(n392), .B(n391), .Z(n404) );
  XOR2_X1 U454 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n394) );
  XNOR2_X1 U455 ( .A(G134GAT), .B(G162GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n402) );
  XOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n396) );
  XNOR2_X1 U458 ( .A(G29GAT), .B(G218GAT), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U460 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n491) );
  NAND2_X1 U467 ( .A1(n409), .A2(n491), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(KEYINPUT47), .ZN(n416) );
  XOR2_X1 U469 ( .A(n518), .B(KEYINPUT76), .Z(n569) );
  INV_X1 U470 ( .A(n584), .ZN(n484) );
  XOR2_X1 U471 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n412) );
  INV_X1 U472 ( .A(n491), .ZN(n573) );
  XNOR2_X1 U473 ( .A(KEYINPUT36), .B(n573), .ZN(n592) );
  NAND2_X1 U474 ( .A1(n588), .A2(n592), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  NAND2_X1 U476 ( .A1(n484), .A2(n413), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n569), .A2(n414), .ZN(n415) );
  NOR2_X1 U478 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT48), .ZN(n560) );
  NOR2_X1 U480 ( .A1(n508), .A2(n560), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n418), .B(KEYINPUT54), .ZN(n440) );
  XOR2_X1 U482 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n420) );
  XNOR2_X1 U483 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n439) );
  XOR2_X1 U485 ( .A(KEYINPUT96), .B(G57GAT), .Z(n424) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U488 ( .A(n425), .B(G85GAT), .Z(n432) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U492 ( .A(G141GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n433), .B(KEYINPUT95), .ZN(n437) );
  XOR2_X1 U495 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n435) );
  XNOR2_X1 U496 ( .A(G162GAT), .B(KEYINPUT92), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n450) );
  XOR2_X1 U498 ( .A(n450), .B(KEYINPUT94), .Z(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n473) );
  XOR2_X1 U501 ( .A(KEYINPUT97), .B(n473), .Z(n533) );
  INV_X1 U502 ( .A(n533), .ZN(n486) );
  NAND2_X1 U503 ( .A1(n440), .A2(n486), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n441), .B(KEYINPUT64), .ZN(n578) );
  XNOR2_X1 U505 ( .A(n442), .B(KEYINPUT81), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n443), .B(G155GAT), .ZN(n447) );
  XOR2_X1 U507 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n445) );
  XNOR2_X1 U508 ( .A(G148GAT), .B(KEYINPUT90), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U510 ( .A(n447), .B(n446), .Z(n457) );
  XOR2_X1 U511 ( .A(G204GAT), .B(KEYINPUT93), .Z(n449) );
  XNOR2_X1 U512 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U514 ( .A(n451), .B(n450), .Z(n453) );
  NAND2_X1 U515 ( .A1(G228GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n476) );
  NOR2_X1 U520 ( .A1(n578), .A2(n476), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT55), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n548), .A2(n574), .ZN(n465) );
  XOR2_X1 U523 ( .A(G176GAT), .B(KEYINPUT56), .Z(n463) );
  XNOR2_X1 U524 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n462) );
  XNOR2_X1 U525 ( .A(KEYINPUT37), .B(KEYINPUT110), .ZN(n483) );
  NOR2_X1 U526 ( .A1(n466), .A2(n476), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT25), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT101), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n476), .A2(n510), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT26), .ZN(n577) );
  XOR2_X1 U531 ( .A(n536), .B(KEYINPUT27), .Z(n477) );
  NOR2_X1 U532 ( .A1(n577), .A2(n477), .ZN(n470) );
  NOR2_X1 U533 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT102), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(KEYINPUT103), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT28), .B(n476), .Z(n514) );
  INV_X1 U538 ( .A(n514), .ZN(n540) );
  OR2_X1 U539 ( .A1(n477), .A2(n486), .ZN(n558) );
  NOR2_X1 U540 ( .A1(n540), .A2(n558), .ZN(n544) );
  NAND2_X1 U541 ( .A1(n544), .A2(n510), .ZN(n478) );
  NAND2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U543 ( .A(KEYINPUT104), .B(n480), .ZN(n494) );
  NAND2_X1 U544 ( .A1(n494), .A2(n592), .ZN(n481) );
  NOR2_X1 U545 ( .A1(n588), .A2(n481), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n532) );
  NAND2_X1 U547 ( .A1(n484), .A2(n569), .ZN(n496) );
  XNOR2_X2 U548 ( .A(n485), .B(KEYINPUT38), .ZN(n515) );
  NOR2_X1 U549 ( .A1(n486), .A2(n515), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n488) );
  INV_X1 U551 ( .A(G29GAT), .ZN(n487) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n498) );
  NAND2_X1 U553 ( .A1(n491), .A2(n588), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT87), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT16), .B(n493), .ZN(n495) );
  NAND2_X1 U556 ( .A1(n495), .A2(n494), .ZN(n519) );
  NOR2_X1 U557 ( .A1(n496), .A2(n519), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n533), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n536), .A2(n504), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT106), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G8GAT), .B(n501), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U565 ( .A1(n504), .A2(n545), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n506) );
  NAND2_X1 U568 ( .A1(n504), .A2(n540), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G22GAT), .B(n507), .ZN(G1327GAT) );
  NOR2_X1 U571 ( .A1(n508), .A2(n515), .ZN(n509) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n509), .Z(G1329GAT) );
  INV_X1 U573 ( .A(KEYINPUT40), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n515), .A2(n510), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n515), .A2(n514), .ZN(n517) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(G1331GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT42), .B(KEYINPUT113), .Z(n521) );
  NAND2_X1 U581 ( .A1(n548), .A2(n518), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n531), .A2(n519), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n527), .A2(n533), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n522), .ZN(G1332GAT) );
  NAND2_X1 U586 ( .A1(n536), .A2(n527), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n525) );
  NAND2_X1 U589 ( .A1(n527), .A2(n545), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT43), .B(KEYINPUT116), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n540), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G78GAT), .B(n530), .ZN(G1335GAT) );
  XOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT117), .Z(n535) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n533), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n541), .A2(n536), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G92GAT), .B(n537), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n541), .A2(n545), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT118), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G99GAT), .B(n539), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U609 ( .A1(n560), .A2(n546), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n569), .A2(n555), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT49), .B(KEYINPUT122), .Z(n550) );
  NAND2_X1 U613 ( .A1(n555), .A2(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT121), .Z(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1341GAT) );
  NAND2_X1 U617 ( .A1(n555), .A2(n571), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT50), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n554), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U621 ( .A1(n555), .A2(n573), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  OR2_X1 U623 ( .A1(n577), .A2(n558), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n566) );
  AND2_X1 U625 ( .A1(n580), .A2(n566), .ZN(n561) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n561), .Z(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U628 ( .A1(n566), .A2(n367), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n588), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U634 ( .A1(n566), .A2(n573), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT58), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(n576), .ZN(G1351GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(n579), .Z(n591) );
  NAND2_X1 U646 ( .A1(n591), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n591), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

