

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772;

  NOR2_X1 U371 ( .A1(n688), .A2(KEYINPUT81), .ZN(n689) );
  XOR2_X1 U372 ( .A(n553), .B(n474), .Z(n349) );
  XOR2_X1 U373 ( .A(n640), .B(KEYINPUT85), .Z(n350) );
  XOR2_X1 U374 ( .A(n628), .B(KEYINPUT82), .Z(n351) );
  XOR2_X1 U375 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n352) );
  XOR2_X1 U376 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n353) );
  AND2_X1 U377 ( .A1(G221), .A2(n540), .ZN(n354) );
  AND2_X2 U378 ( .A1(n427), .A2(n762), .ZN(n688) );
  AND2_X2 U379 ( .A1(n369), .A2(n389), .ZN(n367) );
  OR2_X2 U380 ( .A1(n742), .A2(n371), .ZN(n369) );
  XNOR2_X2 U381 ( .A(n535), .B(n534), .ZN(n697) );
  INV_X1 U382 ( .A(n742), .ZN(n362) );
  XNOR2_X1 U383 ( .A(n373), .B(n350), .ZN(n417) );
  AND2_X1 U384 ( .A1(n372), .A2(KEYINPUT65), .ZN(n364) );
  AND2_X1 U385 ( .A1(n417), .A2(n404), .ZN(n415) );
  AND2_X1 U386 ( .A1(n663), .A2(n358), .ZN(n357) );
  XNOR2_X1 U387 ( .A(n450), .B(n377), .ZN(n485) );
  NOR2_X1 U388 ( .A1(n635), .A2(n399), .ZN(n678) );
  NAND2_X1 U389 ( .A1(n385), .A2(n355), .ZN(n635) );
  NAND2_X1 U390 ( .A1(n693), .A2(n694), .ZN(n589) );
  XNOR2_X1 U391 ( .A(n397), .B(KEYINPUT6), .ZN(n610) );
  XNOR2_X1 U392 ( .A(n384), .B(n349), .ZN(n607) );
  OR2_X1 U393 ( .A1(n730), .A2(G902), .ZN(n457) );
  INV_X1 U394 ( .A(n392), .ZN(n391) );
  NAND2_X1 U395 ( .A1(n650), .A2(n393), .ZN(n392) );
  INV_X1 U396 ( .A(G953), .ZN(n741) );
  INV_X1 U397 ( .A(KEYINPUT3), .ZN(n482) );
  BUF_X1 U398 ( .A(G110), .Z(n440) );
  INV_X1 U399 ( .A(G143), .ZN(n380) );
  INV_X1 U400 ( .A(G125), .ZN(n383) );
  INV_X1 U401 ( .A(KEYINPUT35), .ZN(n377) );
  NAND2_X1 U402 ( .A1(n365), .A2(n364), .ZN(n363) );
  NAND2_X1 U403 ( .A1(n370), .A2(n391), .ZN(n368) );
  NAND2_X1 U404 ( .A1(n416), .A2(n415), .ZN(n370) );
  AND2_X1 U405 ( .A1(n490), .A2(n639), .ZN(n374) );
  OR2_X1 U406 ( .A1(n359), .A2(n351), .ZN(n358) );
  NOR2_X1 U407 ( .A1(n767), .A2(n638), .ZN(n490) );
  XNOR2_X1 U408 ( .A(n485), .B(G122), .ZN(G24) );
  XNOR2_X1 U409 ( .A(n613), .B(KEYINPUT109), .ZN(n767) );
  AND2_X1 U410 ( .A1(n622), .A2(n707), .ZN(n604) );
  NOR2_X1 U411 ( .A1(n463), .A2(n405), .ZN(n462) );
  NOR2_X1 U412 ( .A1(n493), .A2(n491), .ZN(n603) );
  XNOR2_X1 U413 ( .A(n386), .B(n353), .ZN(n385) );
  OR2_X1 U414 ( .A1(n615), .A2(n614), .ZN(n386) );
  XNOR2_X1 U415 ( .A(n382), .B(KEYINPUT106), .ZN(n381) );
  NOR2_X1 U416 ( .A1(n589), .A2(n610), .ZN(n590) );
  NOR2_X1 U417 ( .A1(n610), .A2(n615), .ZN(n382) );
  XNOR2_X1 U418 ( .A(n609), .B(KEYINPUT72), .ZN(n615) );
  NOR2_X1 U419 ( .A1(n607), .A2(n691), .ZN(n694) );
  XOR2_X1 U420 ( .A(n659), .B(n658), .Z(n408) );
  INV_X1 U421 ( .A(n616), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n730), .B(n729), .ZN(n410) );
  XOR2_X1 U423 ( .A(G478), .B(n511), .Z(n623) );
  XNOR2_X1 U424 ( .A(n735), .B(KEYINPUT123), .ZN(n409) );
  OR2_X1 U425 ( .A1(n735), .A2(G902), .ZN(n384) );
  XOR2_X1 U426 ( .A(n661), .B(KEYINPUT62), .Z(n412) );
  XOR2_X1 U427 ( .A(n654), .B(n653), .Z(n411) );
  XOR2_X1 U428 ( .A(n523), .B(n522), .Z(n654) );
  NOR2_X1 U429 ( .A1(n596), .A2(n572), .ZN(n573) );
  NAND2_X1 U430 ( .A1(n390), .A2(KEYINPUT65), .ZN(n389) );
  OR2_X1 U431 ( .A1(n392), .A2(KEYINPUT83), .ZN(n371) );
  INV_X1 U432 ( .A(n650), .ZN(n390) );
  XNOR2_X1 U433 ( .A(n515), .B(n514), .ZN(n521) );
  XNOR2_X1 U434 ( .A(n469), .B(n468), .ZN(n557) );
  XNOR2_X1 U435 ( .A(n564), .B(KEYINPUT10), .ZN(n541) );
  XNOR2_X1 U436 ( .A(n551), .B(KEYINPUT15), .ZN(n648) );
  XNOR2_X1 U437 ( .A(n487), .B(KEYINPUT75), .ZN(n486) );
  XNOR2_X1 U438 ( .A(n482), .B(G116), .ZN(n469) );
  XNOR2_X1 U439 ( .A(n383), .B(G146), .ZN(n564) );
  XNOR2_X1 U440 ( .A(G119), .B(G113), .ZN(n468) );
  XOR2_X1 U441 ( .A(G104), .B(G122), .Z(n513) );
  INV_X1 U442 ( .A(KEYINPUT92), .ZN(n388) );
  INV_X1 U443 ( .A(G953), .ZN(n504) );
  INV_X1 U444 ( .A(KEYINPUT65), .ZN(n393) );
  XNOR2_X2 U445 ( .A(n484), .B(KEYINPUT45), .ZN(n742) );
  NOR2_X2 U446 ( .A1(n398), .A2(n669), .ZN(n471) );
  XNOR2_X2 U447 ( .A(n472), .B(n586), .ZN(n398) );
  NAND2_X1 U448 ( .A1(n356), .A2(n485), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n471), .B(n470), .ZN(n356) );
  NAND2_X2 U450 ( .A1(n360), .A2(n357), .ZN(n484) );
  XNOR2_X1 U451 ( .A(n579), .B(KEYINPUT97), .ZN(n359) );
  XNOR2_X2 U452 ( .A(n361), .B(n591), .ZN(n360) );
  NAND2_X1 U453 ( .A1(n362), .A2(n414), .ZN(n372) );
  NAND2_X2 U454 ( .A1(n366), .A2(n363), .ZN(n652) );
  INV_X1 U455 ( .A(n370), .ZN(n365) );
  AND2_X2 U456 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U457 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X1 U458 ( .A(n637), .B(KEYINPUT46), .ZN(n375) );
  NAND2_X1 U459 ( .A1(n376), .A2(n694), .ZN(n577) );
  NAND2_X1 U460 ( .A1(n387), .A2(n376), .ZN(n453) );
  XNOR2_X1 U461 ( .A(n396), .B(n388), .ZN(n376) );
  XNOR2_X2 U462 ( .A(n378), .B(n499), .ZN(n428) );
  NOR2_X1 U463 ( .A1(n641), .A2(n378), .ZN(n611) );
  NAND2_X2 U464 ( .A1(n592), .A2(n706), .ZN(n378) );
  NAND2_X1 U465 ( .A1(n394), .A2(n473), .ZN(n472) );
  XNOR2_X2 U466 ( .A(n488), .B(n486), .ZN(n394) );
  BUF_X1 U467 ( .A(n669), .Z(n379) );
  XNOR2_X2 U468 ( .A(n380), .B(G128), .ZN(n558) );
  NAND2_X1 U469 ( .A1(n381), .A2(n677), .ZN(n641) );
  INV_X1 U470 ( .A(n607), .ZN(n601) );
  XNOR2_X1 U471 ( .A(n550), .B(n549), .ZN(n735) );
  INV_X1 U472 ( .A(n714), .ZN(n387) );
  NAND2_X1 U473 ( .A1(n394), .A2(n407), .ZN(n464) );
  XNOR2_X1 U474 ( .A(n488), .B(n486), .ZN(n395) );
  XNOR2_X1 U475 ( .A(n575), .B(n574), .ZN(n396) );
  XNOR2_X1 U476 ( .A(n575), .B(n574), .ZN(n466) );
  BUF_X2 U477 ( .A(n697), .Z(n397) );
  BUF_X1 U478 ( .A(n428), .Z(n399) );
  NAND2_X1 U479 ( .A1(n460), .A2(n745), .ZN(n402) );
  NAND2_X1 U480 ( .A1(n400), .A2(n401), .ZN(n403) );
  NAND2_X1 U481 ( .A1(n403), .A2(n402), .ZN(n559) );
  INV_X1 U482 ( .A(n460), .ZN(n400) );
  INV_X1 U483 ( .A(n745), .ZN(n401) );
  XNOR2_X1 U484 ( .A(n526), .B(n525), .ZN(n588) );
  XNOR2_X1 U485 ( .A(n524), .B(G475), .ZN(n525) );
  INV_X1 U486 ( .A(KEYINPUT25), .ZN(n474) );
  XNOR2_X1 U487 ( .A(n538), .B(n539), .ZN(n730) );
  XNOR2_X1 U488 ( .A(n536), .B(n454), .ZN(n498) );
  INV_X1 U489 ( .A(KEYINPUT87), .ZN(n470) );
  XNOR2_X1 U490 ( .A(G902), .B(KEYINPUT89), .ZN(n551) );
  XNOR2_X1 U491 ( .A(KEYINPUT71), .B(G131), .ZN(n532) );
  XOR2_X1 U492 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n518) );
  XNOR2_X1 U493 ( .A(G140), .B(KEYINPUT98), .ZN(n517) );
  NOR2_X1 U494 ( .A1(n770), .A2(n420), .ZN(n419) );
  INV_X1 U495 ( .A(n687), .ZN(n420) );
  XNOR2_X1 U496 ( .A(G119), .B(n440), .ZN(n547) );
  INV_X1 U497 ( .A(KEYINPUT34), .ZN(n452) );
  INV_X1 U498 ( .A(n623), .ZN(n479) );
  NOR2_X1 U499 ( .A1(n587), .A2(KEYINPUT105), .ZN(n463) );
  XNOR2_X1 U500 ( .A(n481), .B(G469), .ZN(n480) );
  INV_X1 U501 ( .A(KEYINPUT74), .ZN(n481) );
  INV_X1 U502 ( .A(G472), .ZN(n534) );
  INV_X1 U503 ( .A(KEYINPUT22), .ZN(n487) );
  INV_X1 U504 ( .A(KEYINPUT44), .ZN(n591) );
  XNOR2_X1 U505 ( .A(n455), .B(G140), .ZN(n542) );
  INV_X1 U506 ( .A(G137), .ZN(n455) );
  OR2_X1 U507 ( .A1(G237), .A2(G902), .ZN(n567) );
  INV_X1 U508 ( .A(KEYINPUT104), .ZN(n423) );
  NOR2_X1 U509 ( .A1(n588), .A2(n623), .ZN(n633) );
  XNOR2_X1 U510 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U511 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n545) );
  XNOR2_X1 U512 ( .A(n544), .B(n543), .ZN(n546) );
  INV_X1 U513 ( .A(KEYINPUT94), .ZN(n543) );
  INV_X1 U514 ( .A(G134), .ZN(n497) );
  INV_X1 U515 ( .A(KEYINPUT83), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n519), .B(n406), .ZN(n520) );
  XNOR2_X1 U517 ( .A(G143), .B(G113), .ZN(n512) );
  XNOR2_X1 U518 ( .A(n542), .B(KEYINPUT93), .ZN(n454) );
  XOR2_X1 U519 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n561) );
  NAND2_X1 U520 ( .A1(n633), .A2(n598), .ZN(n489) );
  XNOR2_X1 U521 ( .A(n504), .B(KEYINPUT64), .ZN(n763) );
  XNOR2_X1 U522 ( .A(n557), .B(n467), .ZN(n746) );
  XNOR2_X1 U523 ( .A(KEYINPUT16), .B(G122), .ZN(n467) );
  INV_X1 U524 ( .A(G107), .ZN(n475) );
  XOR2_X1 U525 ( .A(KEYINPUT102), .B(G107), .Z(n502) );
  XNOR2_X1 U526 ( .A(G116), .B(G122), .ZN(n501) );
  XOR2_X1 U527 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n508) );
  XNOR2_X1 U528 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n456) );
  NAND2_X1 U529 ( .A1(n601), .A2(n492), .ZN(n491) );
  XNOR2_X1 U530 ( .A(n601), .B(KEYINPUT103), .ZN(n690) );
  XNOR2_X1 U531 ( .A(n538), .B(n494), .ZN(n661) );
  XNOR2_X1 U532 ( .A(n496), .B(n495), .ZN(n494) );
  BUF_X1 U533 ( .A(n763), .Z(n445) );
  INV_X1 U534 ( .A(KEYINPUT2), .ZN(n448) );
  NOR2_X1 U535 ( .A1(n722), .A2(n635), .ZN(n636) );
  NOR2_X1 U536 ( .A1(n479), .A2(n626), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n453), .B(n452), .ZN(n451) );
  INV_X1 U538 ( .A(KEYINPUT124), .ZN(n436) );
  INV_X1 U539 ( .A(KEYINPUT60), .ZN(n430) );
  INV_X1 U540 ( .A(KEYINPUT122), .ZN(n434) );
  INV_X1 U541 ( .A(KEYINPUT56), .ZN(n432) );
  AND2_X1 U542 ( .A1(n419), .A2(n413), .ZN(n404) );
  OR2_X1 U543 ( .A1(n601), .A2(n483), .ZN(n405) );
  XOR2_X1 U544 ( .A(n518), .B(n517), .Z(n406) );
  AND2_X1 U545 ( .A1(n587), .A2(KEYINPUT105), .ZN(n407) );
  OR2_X1 U546 ( .A1(n648), .A2(KEYINPUT83), .ZN(n413) );
  NOR2_X1 U547 ( .A1(n445), .A2(G952), .ZN(n738) );
  INV_X1 U548 ( .A(n738), .ZN(n442) );
  NOR2_X1 U549 ( .A1(n395), .A2(KEYINPUT105), .ZN(n465) );
  AND2_X1 U550 ( .A1(n395), .A2(n610), .ZN(n580) );
  AND2_X1 U551 ( .A1(n417), .A2(n419), .ZN(n762) );
  NAND2_X1 U552 ( .A1(n742), .A2(n418), .ZN(n416) );
  AND2_X1 U553 ( .A1(n648), .A2(KEYINPUT83), .ZN(n418) );
  AND2_X1 U554 ( .A1(n421), .A2(n741), .ZN(n449) );
  XNOR2_X1 U555 ( .A(KEYINPUT119), .B(n726), .ZN(n421) );
  NAND2_X1 U556 ( .A1(n697), .A2(KEYINPUT104), .ZN(n424) );
  NAND2_X1 U557 ( .A1(n422), .A2(n423), .ZN(n425) );
  NAND2_X1 U558 ( .A1(n424), .A2(n425), .ZN(n600) );
  INV_X1 U559 ( .A(n697), .ZN(n422) );
  NOR2_X2 U560 ( .A1(n652), .A2(n651), .ZN(n426) );
  BUF_X1 U561 ( .A(n742), .Z(n427) );
  NOR2_X2 U562 ( .A1(n652), .A2(n651), .ZN(n736) );
  BUF_X1 U563 ( .A(n559), .Z(n537) );
  XNOR2_X1 U564 ( .A(n446), .B(KEYINPUT30), .ZN(n493) );
  NOR2_X2 U565 ( .A1(n428), .A2(n573), .ZN(n575) );
  XNOR2_X1 U566 ( .A(n603), .B(n602), .ZN(n622) );
  XNOR2_X1 U567 ( .A(n429), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U568 ( .A1(n438), .A2(n442), .ZN(n429) );
  XNOR2_X1 U569 ( .A(n431), .B(n430), .ZN(G60) );
  NAND2_X1 U570 ( .A1(n439), .A2(n442), .ZN(n431) );
  XNOR2_X1 U571 ( .A(n433), .B(n432), .ZN(G51) );
  NAND2_X1 U572 ( .A1(n441), .A2(n442), .ZN(n433) );
  XNOR2_X1 U573 ( .A(n435), .B(n434), .ZN(G54) );
  NAND2_X1 U574 ( .A1(n444), .A2(n442), .ZN(n435) );
  XNOR2_X1 U575 ( .A(n437), .B(n436), .ZN(G66) );
  NAND2_X1 U576 ( .A1(n443), .A2(n442), .ZN(n437) );
  NAND2_X1 U577 ( .A1(n464), .A2(n462), .ZN(n461) );
  XNOR2_X1 U578 ( .A(n662), .B(n412), .ZN(n438) );
  XNOR2_X1 U579 ( .A(n655), .B(n411), .ZN(n439) );
  XNOR2_X1 U580 ( .A(n737), .B(n409), .ZN(n443) );
  XNOR2_X1 U581 ( .A(n731), .B(n410), .ZN(n444) );
  XNOR2_X1 U582 ( .A(n660), .B(n408), .ZN(n441) );
  NAND2_X1 U583 ( .A1(n600), .A2(n706), .ZN(n446) );
  NAND2_X1 U584 ( .A1(n447), .A2(n725), .ZN(n726) );
  XNOR2_X1 U585 ( .A(n689), .B(n448), .ZN(n447) );
  XNOR2_X1 U586 ( .A(n449), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U587 ( .A1(n451), .A2(n478), .ZN(n450) );
  XNOR2_X2 U588 ( .A(n616), .B(n456), .ZN(n693) );
  XNOR2_X2 U589 ( .A(n457), .B(n480), .ZN(n616) );
  XNOR2_X2 U590 ( .A(n458), .B(n500), .ZN(n592) );
  NAND2_X1 U591 ( .A1(n656), .A2(n566), .ZN(n458) );
  XNOR2_X1 U592 ( .A(n459), .B(n565), .ZN(n656) );
  XNOR2_X1 U593 ( .A(n560), .B(n746), .ZN(n459) );
  XNOR2_X1 U594 ( .A(n460), .B(n529), .ZN(n495) );
  XNOR2_X2 U595 ( .A(n477), .B(KEYINPUT4), .ZN(n460) );
  NOR2_X2 U596 ( .A1(n465), .A2(n461), .ZN(n669) );
  NOR2_X2 U597 ( .A1(n466), .A2(n489), .ZN(n488) );
  NOR2_X1 U598 ( .A1(n702), .A2(n396), .ZN(n576) );
  XNOR2_X1 U599 ( .A(n584), .B(KEYINPUT78), .ZN(n473) );
  XNOR2_X2 U600 ( .A(n476), .B(n475), .ZN(n745) );
  XNOR2_X2 U601 ( .A(G104), .B(G110), .ZN(n476) );
  XNOR2_X2 U602 ( .A(G101), .B(KEYINPUT69), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n498), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n354), .B(n756), .ZN(n550) );
  INV_X1 U605 ( .A(n614), .ZN(n483) );
  NOR2_X1 U606 ( .A1(n616), .A2(n606), .ZN(n492) );
  XNOR2_X1 U607 ( .A(n531), .B(n557), .ZN(n496) );
  XNOR2_X2 U608 ( .A(n754), .B(G146), .ZN(n538) );
  XNOR2_X2 U609 ( .A(n533), .B(n532), .ZN(n754) );
  XNOR2_X2 U610 ( .A(n558), .B(n497), .ZN(n533) );
  BUF_X1 U611 ( .A(n592), .Z(n624) );
  XOR2_X1 U612 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n499) );
  AND2_X1 U613 ( .A1(G210), .A2(n567), .ZN(n500) );
  INV_X1 U614 ( .A(KEYINPUT48), .ZN(n640) );
  XNOR2_X1 U615 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U616 ( .A(KEYINPUT32), .ZN(n585) );
  XNOR2_X1 U617 ( .A(n585), .B(KEYINPUT66), .ZN(n586) );
  XNOR2_X1 U618 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U619 ( .A(n533), .B(n503), .ZN(n510) );
  XOR2_X1 U620 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n506) );
  NAND2_X1 U621 ( .A1(G234), .A2(n763), .ZN(n505) );
  XNOR2_X1 U622 ( .A(n506), .B(n505), .ZN(n540) );
  NAND2_X1 U623 ( .A1(G217), .A2(n540), .ZN(n507) );
  XNOR2_X1 U624 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U625 ( .A(n510), .B(n509), .ZN(n733) );
  NOR2_X1 U626 ( .A1(G902), .A2(n733), .ZN(n511) );
  XNOR2_X1 U627 ( .A(n513), .B(n512), .ZN(n523) );
  NOR2_X1 U628 ( .A1(G953), .A2(G237), .ZN(n530) );
  NAND2_X1 U629 ( .A1(G214), .A2(n530), .ZN(n515) );
  INV_X1 U630 ( .A(n541), .ZN(n514) );
  INV_X1 U631 ( .A(n532), .ZN(n516) );
  XNOR2_X1 U632 ( .A(n516), .B(KEYINPUT12), .ZN(n519) );
  NOR2_X1 U633 ( .A1(G902), .A2(n654), .ZN(n526) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n524) );
  XNOR2_X1 U635 ( .A(KEYINPUT101), .B(n588), .ZN(n527) );
  NAND2_X1 U636 ( .A1(n623), .A2(n527), .ZN(n684) );
  INV_X1 U637 ( .A(n684), .ZN(n671) );
  NOR2_X1 U638 ( .A1(n623), .A2(n527), .ZN(n677) );
  NOR2_X1 U639 ( .A1(n671), .A2(n677), .ZN(n711) );
  INV_X1 U640 ( .A(n711), .ZN(n628) );
  XNOR2_X1 U641 ( .A(G137), .B(KEYINPUT96), .ZN(n528) );
  XNOR2_X1 U642 ( .A(n352), .B(n528), .ZN(n529) );
  NAND2_X1 U643 ( .A1(n530), .A2(G210), .ZN(n531) );
  NOR2_X1 U644 ( .A1(n661), .A2(G902), .ZN(n535) );
  NAND2_X1 U645 ( .A1(G227), .A2(n445), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n541), .B(n542), .ZN(n756) );
  XNOR2_X1 U647 ( .A(G128), .B(KEYINPUT95), .ZN(n544) );
  XNOR2_X1 U648 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U649 ( .A(n648), .ZN(n566) );
  NAND2_X1 U650 ( .A1(G234), .A2(n566), .ZN(n552) );
  XNOR2_X1 U651 ( .A(KEYINPUT20), .B(n552), .ZN(n554) );
  NAND2_X1 U652 ( .A1(G217), .A2(n554), .ZN(n553) );
  NAND2_X1 U653 ( .A1(G221), .A2(n554), .ZN(n555) );
  XOR2_X1 U654 ( .A(KEYINPUT21), .B(n555), .Z(n598) );
  INV_X1 U655 ( .A(n598), .ZN(n691) );
  INV_X1 U656 ( .A(n589), .ZN(n556) );
  NAND2_X1 U657 ( .A1(n397), .A2(n556), .ZN(n702) );
  XNOR2_X1 U658 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U659 ( .A1(G224), .A2(n763), .ZN(n562) );
  XNOR2_X1 U660 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U661 ( .A(n564), .B(n563), .Z(n565) );
  NAND2_X1 U662 ( .A1(G214), .A2(n567), .ZN(n706) );
  NAND2_X1 U663 ( .A1(G234), .A2(G237), .ZN(n568) );
  XNOR2_X1 U664 ( .A(n568), .B(KEYINPUT14), .ZN(n571) );
  NAND2_X1 U665 ( .A1(G952), .A2(n571), .ZN(n569) );
  XNOR2_X1 U666 ( .A(KEYINPUT90), .B(n569), .ZN(n720) );
  NOR2_X1 U667 ( .A1(G953), .A2(n720), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n741), .A2(G898), .ZN(n570) );
  XNOR2_X1 U669 ( .A(n570), .B(KEYINPUT91), .ZN(n751) );
  NAND2_X1 U670 ( .A1(G902), .A2(n571), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n751), .A2(n593), .ZN(n572) );
  INV_X1 U672 ( .A(KEYINPUT0), .ZN(n574) );
  XNOR2_X1 U673 ( .A(n576), .B(KEYINPUT31), .ZN(n683) );
  NOR2_X1 U674 ( .A1(n397), .A2(n577), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n578), .A2(n355), .ZN(n665) );
  NAND2_X1 U676 ( .A1(n683), .A2(n665), .ZN(n579) );
  XOR2_X1 U677 ( .A(KEYINPUT86), .B(n580), .Z(n581) );
  NOR2_X1 U678 ( .A1(n690), .A2(n581), .ZN(n582) );
  INV_X1 U679 ( .A(n693), .ZN(n587) );
  NAND2_X1 U680 ( .A1(n582), .A2(n587), .ZN(n663) );
  NAND2_X1 U681 ( .A1(n690), .A2(n610), .ZN(n583) );
  NOR2_X1 U682 ( .A1(n587), .A2(n583), .ZN(n584) );
  INV_X1 U683 ( .A(n600), .ZN(n614) );
  INV_X1 U684 ( .A(n588), .ZN(n626) );
  XNOR2_X1 U685 ( .A(n590), .B(KEYINPUT33), .ZN(n714) );
  INV_X1 U686 ( .A(n624), .ZN(n646) );
  XNOR2_X1 U687 ( .A(KEYINPUT38), .B(n646), .ZN(n707) );
  OR2_X1 U688 ( .A1(n445), .A2(n593), .ZN(n594) );
  NOR2_X1 U689 ( .A1(G900), .A2(n594), .ZN(n595) );
  NOR2_X1 U690 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U691 ( .A(n597), .B(KEYINPUT79), .ZN(n599) );
  NAND2_X1 U692 ( .A1(n599), .A2(n598), .ZN(n606) );
  INV_X1 U693 ( .A(KEYINPUT77), .ZN(n602) );
  XNOR2_X1 U694 ( .A(n604), .B(KEYINPUT39), .ZN(n631) );
  NOR2_X1 U695 ( .A1(n684), .A2(n631), .ZN(n605) );
  XNOR2_X1 U696 ( .A(KEYINPUT110), .B(n605), .ZN(n770) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(n606), .ZN(n608) );
  NAND2_X1 U698 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U699 ( .A(KEYINPUT36), .B(n611), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n612), .A2(n693), .ZN(n613) );
  INV_X1 U701 ( .A(KEYINPUT47), .ZN(n618) );
  AND2_X1 U702 ( .A1(n628), .A2(n678), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n619), .A2(KEYINPUT82), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n619), .A2(KEYINPUT47), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n621), .A2(n620), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n622), .A2(n627), .ZN(n676) );
  NOR2_X1 U710 ( .A1(KEYINPUT82), .A2(n628), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n678), .A2(n629), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n676), .A2(n630), .ZN(n638) );
  INV_X1 U713 ( .A(n677), .ZN(n681) );
  NOR2_X1 U714 ( .A1(n681), .A2(n631), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(KEYINPUT40), .ZN(n769) );
  INV_X1 U716 ( .A(n633), .ZN(n709) );
  NAND2_X1 U717 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U718 ( .A1(n709), .A2(n710), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n634), .B(KEYINPUT41), .ZN(n722) );
  XNOR2_X1 U720 ( .A(KEYINPUT42), .B(n636), .ZN(n771) );
  NOR2_X1 U721 ( .A1(n769), .A2(n771), .ZN(n637) );
  XNOR2_X1 U722 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n645) );
  INV_X1 U723 ( .A(n641), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n642), .A2(n706), .ZN(n643) );
  NOR2_X1 U725 ( .A1(n693), .A2(n643), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n687) );
  XNOR2_X1 U728 ( .A(KEYINPUT84), .B(n648), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n649), .A2(KEYINPUT2), .ZN(n650) );
  AND2_X1 U730 ( .A1(KEYINPUT2), .A2(n688), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n736), .A2(G475), .ZN(n655) );
  XOR2_X1 U732 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n653) );
  XNOR2_X1 U733 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n659) );
  BUF_X1 U734 ( .A(n656), .Z(n657) );
  XNOR2_X1 U735 ( .A(n657), .B(KEYINPUT54), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n736), .A2(G210), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n736), .A2(G472), .ZN(n662) );
  XNOR2_X1 U738 ( .A(G101), .B(n663), .ZN(G3) );
  NOR2_X1 U739 ( .A1(n681), .A2(n665), .ZN(n664) );
  XOR2_X1 U740 ( .A(G104), .B(n664), .Z(G6) );
  NOR2_X1 U741 ( .A1(n684), .A2(n665), .ZN(n667) );
  XNOR2_X1 U742 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U743 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U744 ( .A(G107), .B(n668), .ZN(G9) );
  XNOR2_X1 U745 ( .A(n379), .B(n440), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n670), .B(KEYINPUT111), .ZN(G12) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U748 ( .A1(n678), .A2(n671), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U750 ( .A(G128), .B(n674), .ZN(G30) );
  XOR2_X1 U751 ( .A(G143), .B(KEYINPUT113), .Z(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(G45) );
  NAND2_X1 U753 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U755 ( .A(G146), .B(n680), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n681), .A2(n683), .ZN(n682) );
  XOR2_X1 U757 ( .A(G113), .B(n682), .Z(G15) );
  NOR2_X1 U758 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U759 ( .A(G116), .B(KEYINPUT115), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n686), .B(n685), .ZN(G18) );
  XNOR2_X1 U761 ( .A(G140), .B(n687), .ZN(G42) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(n692), .Z(n700) );
  XOR2_X1 U764 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n696) );
  OR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n698), .A2(n397), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(KEYINPUT51), .B(n703), .ZN(n704) );
  NOR2_X1 U771 ( .A1(n722), .A2(n704), .ZN(n705) );
  XOR2_X1 U772 ( .A(KEYINPUT117), .B(n705), .Z(n717) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n715) );
  NOR2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U779 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n721), .B(KEYINPUT118), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n722), .A2(n714), .ZN(n723) );
  NOR2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U784 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n728) );
  XNOR2_X1 U785 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n727) );
  XNOR2_X1 U786 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U787 ( .A1(n426), .A2(G469), .ZN(n731) );
  NAND2_X1 U788 ( .A1(G478), .A2(n426), .ZN(n732) );
  XNOR2_X1 U789 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U790 ( .A1(n738), .A2(n734), .ZN(G63) );
  NAND2_X1 U791 ( .A1(n426), .A2(G217), .ZN(n737) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n740), .A2(G898), .ZN(n744) );
  NAND2_X1 U795 ( .A1(n427), .A2(n741), .ZN(n743) );
  NAND2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n753) );
  BUF_X1 U797 ( .A(n745), .Z(n749) );
  XNOR2_X1 U798 ( .A(G101), .B(n746), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n747), .B(KEYINPUT125), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U802 ( .A(n753), .B(n752), .Z(G69) );
  XOR2_X1 U803 ( .A(n754), .B(KEYINPUT4), .Z(n755) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n761) );
  INV_X1 U805 ( .A(n761), .ZN(n757) );
  XNOR2_X1 U806 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G900), .ZN(n759) );
  XNOR2_X1 U808 ( .A(KEYINPUT126), .B(n759), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n760), .A2(G953), .ZN(n766) );
  XNOR2_X1 U810 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(n445), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U813 ( .A(G125), .B(n767), .ZN(n768) );
  XNOR2_X1 U814 ( .A(n768), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U815 ( .A(n398), .B(G119), .Z(G21) );
  XOR2_X1 U816 ( .A(n769), .B(G131), .Z(G33) );
  XOR2_X1 U817 ( .A(G134), .B(n770), .Z(G36) );
  XNOR2_X1 U818 ( .A(G137), .B(KEYINPUT127), .ZN(n772) );
  XNOR2_X1 U819 ( .A(n772), .B(n771), .ZN(G39) );
endmodule

