//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G140), .Z(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT10), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT65), .A2(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT65), .A2(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(new_n196), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT83), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT65), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(G143), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G146), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n199), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(new_n194), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n204), .B(new_n208), .C1(new_n211), .C2(new_n193), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n209), .A3(G128), .A4(new_n199), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n202), .A2(KEYINPUT82), .A3(new_n209), .A4(G128), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n203), .A2(new_n212), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n221));
  OAI211_X1 g035(.A(G104), .B(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G107), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n224), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n223), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n217), .A2(KEYINPUT84), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT84), .B1(new_n217), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n192), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT11), .B1(new_n236), .B2(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G137), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT11), .A2(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n194), .A2(G143), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n210), .B2(new_n194), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n193), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  INV_X1    g069(.A(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n197), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n253), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n213), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n232), .ZN(new_n261));
  INV_X1    g075(.A(new_n221), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n228), .B1(new_n262), .B2(new_n219), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n226), .A2(new_n225), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT81), .B(G101), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n227), .A3(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(KEYINPUT81), .A3(new_n268), .A4(G101), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT0), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(new_n193), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n270), .A2(new_n193), .A3(KEYINPUT64), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n197), .B2(new_n256), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n273), .B2(new_n202), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT64), .B1(new_n270), .B2(new_n193), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n266), .A2(new_n269), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n261), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n235), .A2(new_n250), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n260), .A2(new_n232), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n233), .B2(new_n234), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n282), .A2(KEYINPUT12), .A3(new_n249), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n282), .B2(new_n249), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n191), .B(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n217), .A2(new_n232), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT84), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n217), .A2(KEYINPUT84), .A3(new_n232), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n280), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n292), .B2(new_n250), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n282), .A2(KEYINPUT12), .A3(new_n249), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n191), .B1(new_n295), .B2(new_n279), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n190), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n250), .A2(KEYINPUT86), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n235), .A2(new_n278), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n235), .B2(new_n278), .ZN(new_n300));
  OR3_X1    g114(.A1(new_n299), .A2(new_n300), .A3(new_n190), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(G469), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n190), .B1(new_n299), .B2(new_n300), .ZN(new_n305));
  INV_X1    g119(.A(new_n190), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(KEYINPUT87), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n279), .A2(new_n306), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n295), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n303), .B(new_n304), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(G469), .A2(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G210), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G224), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AND4_X1   g133(.A1(new_n209), .A2(new_n207), .A3(G128), .A4(new_n199), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT68), .B1(new_n252), .B2(new_n253), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n257), .A2(new_n258), .A3(new_n255), .ZN(new_n322));
  AOI211_X1 g136(.A(G125), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n274), .B2(new_n276), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n323), .A2(KEYINPUT88), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n274), .A2(new_n276), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G125), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n324), .B(new_n213), .C1(new_n254), .C2(new_n259), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n319), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT88), .B1(new_n323), .B2(new_n325), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n327), .A3(new_n330), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n318), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G116), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G119), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G116), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(KEYINPUT69), .A3(G119), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT2), .B(G113), .Z(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n266), .A2(new_n269), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(KEYINPUT5), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(G113), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n343), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n230), .A4(new_n227), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n351), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n332), .A2(new_n335), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n304), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n318), .B1(KEYINPUT89), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(KEYINPUT89), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n323), .B2(new_n325), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n330), .A4(new_n319), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n348), .A2(G113), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n342), .B2(KEYINPUT5), .ZN(new_n368));
  INV_X1    g182(.A(new_n350), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n231), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n351), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n353), .B(KEYINPUT8), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n365), .A2(new_n366), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n356), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n329), .A2(new_n330), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n377), .A2(new_n364), .B1(new_n371), .B2(new_n372), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n374), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n316), .B1(new_n361), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n365), .A2(new_n366), .A3(new_n373), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT90), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n356), .A3(new_n375), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n384), .A2(new_n304), .A3(new_n360), .A4(new_n315), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G214), .B1(G237), .B2(G902), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  OAI21_X1  g204(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n314), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G472), .A2(G902), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G134), .B1(new_n240), .B2(new_n242), .ZN(new_n395));
  INV_X1    g209(.A(new_n238), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n248), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n260), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n249), .A2(new_n274), .A3(new_n276), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n321), .A2(new_n322), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n403), .B2(new_n213), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n249), .A2(new_n274), .A3(KEYINPUT67), .A4(new_n276), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n344), .B(new_n402), .C1(new_n408), .C2(KEYINPUT30), .ZN(new_n409));
  INV_X1    g223(.A(new_n344), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n401), .B(new_n410), .C1(new_n411), .C2(new_n398), .ZN(new_n412));
  INV_X1    g226(.A(G237), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n187), .A2(G210), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT26), .B(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n416), .A2(new_n417), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n409), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n409), .A2(KEYINPUT31), .A3(new_n412), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT71), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n419), .B2(new_n420), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n414), .B(KEYINPUT27), .ZN(new_n429));
  INV_X1    g243(.A(new_n417), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n431), .A3(KEYINPUT71), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n406), .A2(new_n407), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n344), .B1(new_n434), .B2(new_n404), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n400), .A2(new_n437), .A3(new_n410), .A4(new_n401), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n433), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n394), .B1(new_n426), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n418), .A2(new_n431), .A3(KEYINPUT29), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n401), .B1(new_n411), .B2(new_n398), .ZN(new_n444));
  AOI221_X4 g258(.A(new_n443), .B1(new_n344), .B2(new_n444), .C1(new_n436), .C2(new_n438), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT73), .B1(new_n445), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n344), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n447), .B(new_n304), .C1(new_n449), .C2(new_n443), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n421), .B1(new_n409), .B2(new_n412), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n435), .A2(new_n433), .A3(new_n439), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT29), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n446), .B(new_n450), .C1(new_n451), .C2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n442), .A2(KEYINPUT32), .B1(G472), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n440), .B1(new_n424), .B2(new_n425), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n394), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT72), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n457), .C1(new_n458), .C2(new_n394), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G217), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(G234), .B2(new_n304), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT25), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G137), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G140), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT16), .ZN(new_n473));
  XNOR2_X1  g287(.A(G125), .B(G140), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(KEYINPUT16), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n194), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n193), .A2(G119), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(KEYINPUT74), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT74), .B1(new_n339), .B2(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n339), .A2(G128), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(KEYINPUT23), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT75), .B(G110), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n480), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT24), .B(G110), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n486), .A2(KEYINPUT76), .A3(new_n489), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n478), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n475), .B(new_n194), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n487), .A2(new_n488), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n481), .A2(new_n484), .ZN(new_n498));
  INV_X1    g312(.A(G110), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT77), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n496), .A2(new_n500), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n503), .A2(new_n494), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n470), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(new_n501), .A3(KEYINPUT77), .ZN(new_n507));
  INV_X1    g321(.A(new_n470), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n467), .B1(new_n510), .B2(G902), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n504), .B1(new_n503), .B2(new_n494), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n505), .A2(new_n470), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT25), .A3(new_n304), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n466), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n466), .A2(new_n304), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT78), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n509), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n463), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  INV_X1    g341(.A(G953), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT70), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G953), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n529), .A2(new_n531), .A3(G214), .A4(new_n413), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n201), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT91), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n187), .A2(G143), .A3(G214), .A4(new_n413), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n536), .A3(new_n201), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT18), .A2(G131), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n534), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n474), .B(new_n194), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n535), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n536), .B1(new_n532), .B2(new_n201), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n539), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT94), .B(G104), .Z(new_n546));
  XNOR2_X1  g360(.A(G113), .B(G122), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n534), .A2(new_n247), .A3(new_n535), .A4(new_n537), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n543), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n496), .B1(new_n543), .B2(new_n549), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n545), .B(new_n548), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n550), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n475), .A2(G146), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n324), .A2(G140), .ZN(new_n557));
  AND2_X1   g371(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n558));
  NOR2_X1   g372(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n472), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT19), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(KEYINPUT93), .C1(new_n561), .C2(new_n474), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(KEYINPUT93), .B2(new_n560), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n556), .B1(new_n563), .B2(new_n194), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n555), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n548), .B1(new_n565), .B2(new_n545), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n527), .B1(new_n554), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n545), .ZN(new_n568));
  INV_X1    g382(.A(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT95), .A3(new_n553), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n526), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n554), .A2(new_n566), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n526), .A2(KEYINPUT20), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n545), .B1(new_n551), .B2(new_n552), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n569), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n579), .B2(new_n553), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT96), .B(G475), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n390), .A2(new_n464), .A3(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n201), .A2(G128), .ZN(new_n587));
  INV_X1    g401(.A(G134), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n193), .A2(G143), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G122), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT97), .B1(new_n591), .B2(G116), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n336), .A3(G122), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(G116), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n595), .A2(new_n218), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n218), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n590), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n589), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n210), .A2(new_n193), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(KEYINPUT13), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n587), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n587), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n599), .B1(new_n608), .B2(G134), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n601), .A2(G134), .A3(new_n600), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n595), .A2(KEYINPUT14), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n595), .A2(KEYINPUT14), .B1(G116), .B2(new_n591), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n218), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n612), .A2(new_n615), .A3(new_n597), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n586), .B1(new_n609), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G134), .B1(new_n601), .B2(new_n600), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n597), .B1(new_n618), .B2(new_n590), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n613), .A2(new_n614), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n218), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n601), .B2(KEYINPUT13), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n605), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n588), .B1(new_n623), .B2(new_n602), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n621), .B(new_n585), .C1(new_n624), .C2(new_n599), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n617), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n628), .B(G902), .C1(new_n617), .C2(new_n625), .ZN(new_n629));
  INV_X1    g443(.A(G478), .ZN(new_n630));
  OAI22_X1  g444(.A1(new_n627), .A2(new_n629), .B1(KEYINPUT15), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(KEYINPUT15), .ZN(new_n632));
  INV_X1    g446(.A(new_n626), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n628), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n187), .ZN(new_n636));
  NAND2_X1  g450(.A1(G234), .A2(G237), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(G902), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT21), .B(G898), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n637), .A2(G952), .A3(new_n528), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n584), .A2(new_n635), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n392), .A2(new_n524), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G101), .ZN(G3));
  AND2_X1   g461(.A1(new_n314), .A2(new_n391), .ZN(new_n648));
  INV_X1    g462(.A(new_n442), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n458), .B2(G902), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n523), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n617), .A2(new_n625), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT33), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(KEYINPUT33), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(G478), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n630), .A2(new_n304), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n626), .B2(new_n630), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n584), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n662), .A2(new_n388), .A3(new_n644), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n653), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND2_X1  g480(.A1(new_n635), .A2(new_n583), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n643), .B(KEYINPUT103), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n326), .A2(new_n331), .A3(new_n319), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n318), .B1(new_n333), .B2(new_n334), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n357), .A2(new_n359), .ZN(new_n672));
  AOI21_X1  g486(.A(G902), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n315), .B1(new_n673), .B2(new_n384), .ZN(new_n674));
  INV_X1    g488(.A(new_n385), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n387), .B(new_n668), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n572), .B2(new_n573), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n570), .A2(KEYINPUT95), .A3(new_n553), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT95), .B1(new_n570), .B2(new_n553), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n525), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n575), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n678), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT102), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n682), .A3(new_n686), .A4(new_n683), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n667), .B(new_n676), .C1(new_n685), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n653), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT35), .B(G107), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  NAND4_X1  g505(.A1(new_n314), .A2(new_n645), .A3(new_n389), .A4(new_n391), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n649), .A2(new_n650), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT25), .B1(new_n515), .B2(new_n304), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n513), .A2(new_n514), .A3(new_n467), .A4(G902), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n465), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n495), .A2(new_n501), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n508), .A2(KEYINPUT36), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n519), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n692), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT37), .B(G110), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT104), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G12));
  NAND2_X1  g521(.A1(new_n463), .A2(new_n702), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n392), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n685), .A2(new_n687), .ZN(new_n711));
  INV_X1    g525(.A(new_n667), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n641), .B1(new_n638), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n193), .ZN(G30));
  INV_X1    g532(.A(new_n387), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n631), .B2(new_n634), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n584), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n386), .B(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n702), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n714), .B(KEYINPUT39), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n648), .A2(new_n726), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n721), .B(new_n725), .C1(new_n727), .C2(KEYINPUT40), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n448), .A2(new_n412), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n422), .B1(new_n433), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n304), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n442), .A2(KEYINPUT32), .B1(G472), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n460), .A3(new_n462), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n728), .B(new_n734), .C1(KEYINPUT40), .C2(new_n727), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n210), .B(KEYINPUT107), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G45));
  NAND3_X1  g551(.A1(new_n584), .A2(new_n661), .A3(new_n715), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n710), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n194), .ZN(G48));
  OAI21_X1  g554(.A(new_n304), .B1(new_n308), .B2(new_n311), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n391), .A3(new_n312), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n463), .A3(new_n523), .A4(new_n663), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n688), .A2(new_n743), .A3(new_n463), .A4(new_n523), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  AND4_X1   g562(.A1(new_n389), .A2(new_n742), .A3(new_n391), .A4(new_n312), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n463), .A3(new_n645), .A4(new_n702), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NOR2_X1   g565(.A1(new_n574), .A2(new_n576), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n681), .B2(KEYINPUT20), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n386), .B(new_n720), .C1(new_n753), .C2(new_n582), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n584), .A2(KEYINPUT108), .A3(new_n386), .A4(new_n720), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n433), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n449), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n426), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n393), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n523), .A2(new_n762), .A3(new_n650), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n743), .A2(new_n758), .A3(new_n668), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND3_X1  g579(.A1(new_n702), .A2(new_n762), .A3(new_n650), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n738), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n389), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n742), .A2(new_n389), .A3(new_n391), .A4(new_n312), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n762), .A2(new_n650), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n660), .B(new_n714), .C1(new_n577), .C2(new_n583), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n702), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  NOR2_X1   g590(.A1(new_n386), .A2(new_n719), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n391), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n313), .B(KEYINPUT110), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n312), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n297), .A2(KEYINPUT111), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n190), .C1(new_n286), .C2(new_n296), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(G469), .A3(new_n301), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n778), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n785), .A2(new_n524), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n426), .A2(new_n441), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n393), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n455), .A2(G472), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n459), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n772), .A3(new_n523), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n788), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NAND2_X1  g610(.A1(new_n716), .A2(KEYINPUT112), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n711), .A2(new_n798), .A3(new_n712), .A4(new_n715), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n524), .A3(new_n785), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  AND4_X1   g615(.A1(KEYINPUT45), .A2(new_n781), .A3(new_n301), .A4(new_n783), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n297), .B2(new_n301), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n802), .A2(new_n303), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n779), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT46), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n312), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n391), .A3(new_n726), .ZN(new_n812));
  INV_X1    g626(.A(new_n777), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n577), .A2(new_n583), .A3(new_n661), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT43), .Z(new_n817));
  OR3_X1    g631(.A1(new_n817), .A2(new_n694), .A3(new_n724), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n236), .ZN(G39));
  NOR4_X1   g637(.A1(new_n463), .A2(new_n523), .A3(new_n813), .A4(new_n738), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT114), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n391), .B1(new_n809), .B2(new_n810), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT47), .B(new_n391), .C1(new_n809), .C2(new_n810), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n471), .ZN(G42));
  AND2_X1   g646(.A1(new_n742), .A2(new_n312), .ZN(new_n833));
  INV_X1    g647(.A(new_n391), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n771), .A2(new_n523), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n817), .A2(new_n642), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n777), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n743), .A2(new_n777), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT119), .Z(new_n843));
  NOR2_X1   g657(.A1(new_n817), .A2(new_n642), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n702), .A3(new_n771), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT120), .Z(new_n846));
  NOR2_X1   g660(.A1(new_n723), .A2(new_n387), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n743), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT50), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n734), .A2(new_n517), .A3(new_n522), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n641), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n577), .A2(new_n583), .A3(new_n660), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n839), .B2(new_n840), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT51), .B1(new_n841), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n528), .A2(G952), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n838), .B2(new_n749), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n843), .A2(new_n844), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n792), .A2(new_n523), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(new_n865));
  OAI221_X1 g679(.A(new_n859), .B1(new_n662), .B2(new_n851), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n846), .A2(new_n854), .A3(KEYINPUT51), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n867), .B2(new_n839), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  INV_X1    g683(.A(new_n645), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n770), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n742), .A2(new_n391), .A3(new_n312), .A4(new_n668), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n837), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n709), .A2(new_n871), .B1(new_n873), .B2(new_n758), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(KEYINPUT115), .A3(new_n744), .A4(new_n747), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n750), .A2(new_n747), .A3(new_n744), .A4(new_n764), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n577), .A2(new_n583), .A3(new_n635), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n676), .B1(new_n662), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n314), .A3(new_n651), .A4(new_n391), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n463), .A2(new_n523), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n692), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n704), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n635), .A2(new_n714), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n777), .A2(new_n583), .A3(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n391), .A2(new_n887), .A3(new_n314), .A4(new_n711), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n709), .B1(new_n767), .B2(new_n785), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n795), .A2(new_n800), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n716), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n392), .B(new_n709), .C1(new_n892), .C2(new_n772), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n780), .A2(new_n784), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n702), .A2(new_n834), .A3(new_n714), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n733), .A3(new_n758), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n775), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n869), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n901), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n778), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n894), .A2(new_n793), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n785), .A2(new_n524), .A3(new_n786), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n910), .A2(new_n889), .A3(new_n911), .A4(new_n800), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n885), .A3(new_n878), .A4(new_n875), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT53), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n900), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n897), .B(KEYINPUT52), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n869), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n876), .A2(new_n869), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n800), .A2(new_n910), .A3(new_n911), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n885), .A4(new_n889), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n907), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n868), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  OAI22_X1  g740(.A1(new_n857), .A2(new_n926), .B1(G952), .B2(G953), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT49), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n833), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n833), .A2(new_n928), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n723), .A2(new_n719), .A3(new_n814), .A4(new_n834), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n850), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n187), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n891), .B2(new_n899), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n921), .B1(new_n906), .B2(new_n905), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n304), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n671), .A2(new_n672), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n360), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n935), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n940), .B2(new_n945), .ZN(G51));
  OAI21_X1  g761(.A(KEYINPUT54), .B1(new_n936), .B2(new_n937), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(KEYINPUT122), .A3(new_n925), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(KEYINPUT54), .C1(new_n936), .C2(new_n937), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n779), .B(KEYINPUT57), .Z(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n308), .A2(new_n311), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n939), .A2(new_n804), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n953), .A2(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n934), .B1(new_n958), .B2(new_n960), .ZN(G54));
  NAND3_X1  g775(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n679), .A2(new_n680), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n934), .ZN(G60));
  AND2_X1   g780(.A1(new_n655), .A2(new_n656), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n916), .A2(new_n925), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n658), .B(KEYINPUT59), .Z(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n968), .A2(new_n949), .A3(new_n951), .A4(new_n970), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n934), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n938), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n700), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n977), .B(new_n935), .C1(new_n515), .C2(new_n976), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g793(.A(G953), .B1(new_n639), .B2(new_n317), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT124), .ZN(new_n981));
  INV_X1    g795(.A(new_n879), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n885), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n983), .B2(new_n187), .ZN(new_n984));
  INV_X1    g798(.A(new_n672), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(G898), .B2(new_n187), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n984), .B(new_n987), .ZN(G69));
  AOI21_X1  g802(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT126), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n822), .A2(new_n831), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n893), .A2(new_n775), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n920), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n812), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n862), .B1(new_n756), .B2(new_n757), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n402), .B1(new_n408), .B2(KEYINPUT30), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n563), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n187), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI22_X1  g816(.A1(new_n998), .A2(new_n1002), .B1(new_n713), .B2(new_n636), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n662), .A2(new_n880), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n727), .A2(new_n883), .A3(new_n813), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n735), .A2(new_n993), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n636), .B1(new_n992), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(new_n1000), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n991), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1003), .B(new_n990), .C1(new_n1000), .C2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(new_n409), .A2(new_n412), .ZN(new_n1016));
  INV_X1    g830(.A(new_n983), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n992), .A2(new_n997), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  AOI211_X1 g834(.A(new_n421), .B(new_n1016), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1016), .A2(new_n421), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n992), .A2(new_n1010), .A3(new_n1017), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n1020), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1016), .A2(new_n419), .A3(new_n420), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1020), .B1(new_n1025), .B2(new_n451), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT127), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n915), .A2(new_n1027), .ZN(new_n1028));
  NOR4_X1   g842(.A1(new_n1021), .A2(new_n934), .A3(new_n1024), .A4(new_n1028), .ZN(G57));
endmodule


