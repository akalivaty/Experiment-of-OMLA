//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n466));
  XOR2_X1   g041(.A(new_n466), .B(KEYINPUT67), .Z(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(G137), .A3(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n461), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n484), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n462), .A2(G138), .A3(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n491), .A2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n496), .A3(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(G88), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n504), .A2(new_n505), .B1(G50), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n499), .A2(new_n501), .ZN(new_n514));
  INV_X1    g089(.A(new_n497), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n512), .A2(new_n519), .A3(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n502), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n502), .A2(new_n503), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT72), .A4(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n532), .B1(new_n537), .B2(G51), .ZN(G168));
  AOI22_X1  g113(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n534), .A2(G52), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n502), .A2(G90), .A3(new_n503), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n502), .B2(G56), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI211_X1 g126(.A(KEYINPUT74), .B(new_n548), .C1(new_n502), .C2(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n514), .A2(G56), .A3(new_n515), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT74), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(new_n550), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .A4(G651), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n537), .A2(G43), .B1(new_n504), .B2(G81), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G860), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n510), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n503), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n531), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n502), .A2(G65), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n506), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n504), .A2(G91), .B1(new_n569), .B2(new_n571), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n579), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G168), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  OAI21_X1  g163(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n511), .A2(G49), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n531), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n511), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n502), .A2(G86), .A3(new_n503), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n506), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n537), .A2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n504), .A2(G85), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n506), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n537), .B2(G54), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n531), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  AOI21_X1  g200(.A(new_n618), .B1(G559), .B2(new_n560), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT81), .ZN(G148));
  OR2_X1    g202(.A1(new_n618), .A2(G559), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(new_n559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(G868), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g207(.A1(G123), .A2(new_n478), .B1(new_n475), .B2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n634), .A2(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n635), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n654), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT84), .Z(G401));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n444), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT17), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n670), .B1(new_n668), .B2(KEYINPUT85), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(KEYINPUT85), .B2(new_n668), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n671), .B(new_n670), .C1(new_n444), .C2(new_n667), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n640), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n645), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  AND2_X1   g277(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n703));
  NOR2_X1   g278(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT90), .B(G16), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(G166), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G22), .B2(new_n708), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(G1971), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(G1971), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT92), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(KEYINPUT92), .A3(new_n712), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G23), .ZN(new_n717));
  INV_X1    g292(.A(G288), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n716), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT33), .Z(new_n720));
  INV_X1    g295(.A(G1976), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n714), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n601), .A2(G16), .A3(new_n602), .ZN(new_n724));
  OR2_X1    g299(.A1(G6), .A2(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT32), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n724), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G1981), .ZN(new_n731));
  INV_X1    g306(.A(G1981), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n727), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT93), .B1(new_n723), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n715), .A2(new_n722), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n713), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(new_n733), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(KEYINPUT34), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G24), .B(G290), .S(new_n708), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G1986), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G1986), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G25), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n475), .A2(G131), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n478), .A2(G119), .ZN(new_n749));
  NOR2_X1   g324(.A1(G95), .A2(G2105), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT89), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n744), .A2(new_n745), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n741), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT34), .ZN(new_n761));
  INV_X1    g336(.A(new_n740), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n706), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n764), .A2(new_n741), .A3(new_n758), .A4(new_n703), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n767));
  INV_X1    g342(.A(G129), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n477), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  AOI211_X1 g347(.A(new_n769), .B(new_n772), .C1(G141), .C2(new_n475), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(new_n746), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n746), .B2(G32), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT31), .B(G11), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n639), .A2(new_n746), .ZN(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT30), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT102), .Z(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n778), .B(new_n779), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n746), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n786), .B(new_n787), .Z(new_n788));
  INV_X1    g363(.A(G128), .ZN(new_n789));
  INV_X1    g364(.A(G140), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n789), .A2(new_n477), .B1(new_n474), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n794));
  OAI221_X1 g369(.A(G2104), .B1(G116), .B2(new_n464), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n788), .B1(G29), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n775), .A2(new_n776), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n777), .A2(new_n784), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n619), .A2(new_n716), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G4), .B2(new_n716), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT95), .B(G1348), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT100), .B(KEYINPUT24), .ZN(new_n807));
  AOI21_X1  g382(.A(G29), .B1(new_n807), .B2(G34), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G34), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G160), .B2(new_n746), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2084), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n746), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n746), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  NAND2_X1  g390(.A1(G164), .A2(G29), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G27), .B2(G29), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n815), .A2(G2090), .B1(new_n443), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n716), .A2(G21), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G168), .B2(new_n716), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1966), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n746), .A2(G33), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT25), .Z(new_n825));
  INV_X1    g400(.A(G139), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n474), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n462), .A2(G127), .ZN(new_n828));
  AND2_X1   g403(.A1(G115), .A2(G2104), .ZN(new_n829));
  OAI21_X1  g404(.A(G2105), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n823), .B1(new_n833), .B2(G29), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n442), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n815), .B2(G2090), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n834), .A2(new_n442), .B1(new_n817), .B2(new_n443), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n805), .A2(new_n812), .A3(new_n822), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n716), .A2(G5), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G171), .B2(new_n716), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1961), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n708), .A2(G19), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n630), .B2(new_n708), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1341), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n707), .A2(G20), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT23), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n623), .B2(new_n716), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1956), .ZN(new_n849));
  NOR4_X1   g424(.A1(new_n839), .A2(new_n842), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n766), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n765), .A2(new_n851), .ZN(G311));
  INV_X1    g427(.A(new_n764), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n705), .B1(new_n853), .B2(new_n759), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n766), .A3(new_n850), .ZN(G150));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT103), .B(G93), .Z(new_n857));
  OAI22_X1  g432(.A1(new_n536), .A2(new_n856), .B1(new_n531), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n506), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n559), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n553), .A2(new_n861), .A3(new_n557), .A4(new_n558), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n619), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT104), .ZN(new_n871));
  AOI21_X1  g446(.A(G860), .B1(new_n868), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n862), .A2(G860), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  XOR2_X1   g456(.A(G164), .B(new_n797), .Z(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n833), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n882), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n478), .A2(G130), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT108), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n475), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(new_n643), .Z(new_n892));
  OR2_X1    g467(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n753), .B(new_n773), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n896), .A3(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(KEYINPUT106), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n482), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n639), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT109), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n898), .A2(new_n906), .A3(new_n903), .A4(new_n899), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n900), .B2(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g486(.A(G868), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n862), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n618), .B1(new_n579), .B2(new_n585), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n578), .A2(new_n612), .A3(new_n584), .A4(new_n617), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(new_n915), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n578), .A2(new_n584), .B1(new_n612), .B2(new_n617), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n865), .B(new_n628), .Z(new_n923));
  MUX2_X1   g498(.A(new_n916), .B(new_n922), .S(new_n923), .Z(new_n924));
  NOR2_X1   g499(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G166), .B(new_n718), .ZN(new_n927));
  NAND2_X1  g502(.A1(G290), .A2(KEYINPUT110), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n605), .A2(new_n606), .A3(new_n929), .A4(new_n607), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n601), .A2(new_n931), .A3(new_n602), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n602), .B2(new_n601), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(G305), .A2(new_n928), .A3(new_n930), .ZN(new_n936));
  XNOR2_X1  g511(.A(G166), .B(G288), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(KEYINPUT111), .B2(KEYINPUT42), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n926), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n913), .B1(new_n941), .B2(new_n912), .ZN(G295));
  OAI21_X1  g517(.A(new_n913), .B1(new_n941), .B2(new_n912), .ZN(G331));
  OAI211_X1 g518(.A(KEYINPUT112), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(G168), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n541), .A2(new_n542), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT73), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n542), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT112), .B1(new_n950), .B2(new_n540), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(G171), .A2(KEYINPUT112), .A3(G168), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n865), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g530(.A1(G301), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(G168), .A3(new_n944), .ZN(new_n957));
  NAND3_X1  g532(.A1(G286), .A2(new_n955), .A3(G301), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n863), .A3(new_n864), .A4(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n916), .A3(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n954), .A2(new_n959), .B1(new_n920), .B2(new_n921), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n939), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(new_n939), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n961), .B2(new_n960), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT113), .B1(new_n960), .B2(new_n961), .ZN(new_n968));
  INV_X1    g543(.A(new_n959), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n957), .A2(new_n958), .B1(new_n863), .B2(new_n864), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n922), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n954), .A2(new_n916), .A3(new_n959), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n965), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n963), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n964), .B1(new_n975), .B2(new_n963), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT114), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT44), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n964), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT115), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n989));
  INV_X1    g564(.A(new_n981), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n963), .A2(new_n966), .A3(new_n964), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n980), .B2(KEYINPUT114), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n988), .B(new_n989), .C1(new_n993), .C2(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT62), .ZN(new_n996));
  INV_X1    g571(.A(new_n465), .ZN(new_n997));
  INV_X1    g572(.A(new_n472), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT68), .B1(new_n467), .B2(new_n468), .ZN(new_n999));
  OAI211_X1 g574(.A(G40), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n491), .B2(new_n494), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G2084), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1000), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n488), .A2(new_n490), .ZN(new_n1010));
  INV_X1    g585(.A(new_n494), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1966), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(G286), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1000), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(G168), .A3(new_n1006), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1015), .A2(new_n1021), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n996), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT123), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT62), .A3(new_n1027), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1003), .A2(new_n1034), .A3(new_n1005), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1971), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n522), .A2(G8), .A3(new_n523), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1018), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1041), .A2(G1971), .B1(new_n1042), .B2(G2090), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1038), .B(KEYINPUT55), .Z(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(G8), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n595), .A2(G651), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n511), .A2(G48), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1048), .B2(new_n597), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n596), .A2(new_n598), .A3(new_n732), .A4(new_n599), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1012), .A2(G160), .A3(G40), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n718), .A2(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n721), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(G8), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(G8), .B(new_n1060), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT116), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1057), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1040), .A2(new_n1045), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT124), .B1(new_n1018), .B2(G2078), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT53), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT124), .B(new_n1073), .C1(new_n1018), .C2(G2078), .ZN(new_n1074));
  INV_X1    g649(.A(G1961), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1042), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1030), .A2(new_n1033), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n718), .A2(new_n721), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1050), .B1(new_n1058), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1084), .A2(new_n1085), .B1(new_n1087), .B2(new_n1055), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1044), .B1(new_n1043), .B2(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1020), .A2(new_n1006), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G286), .A2(new_n1054), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1067), .A2(new_n1090), .A3(new_n1057), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT63), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(KEYINPUT63), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1070), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1083), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(new_n1066), .A3(new_n1069), .A4(new_n1096), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT117), .A3(new_n1093), .A4(new_n1088), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1030), .A2(new_n1033), .A3(KEYINPUT125), .A4(new_n1079), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n580), .A2(new_n582), .B1(KEYINPUT119), .B2(KEYINPUT57), .ZN(new_n1105));
  NOR2_X1   g680(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT120), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1105), .B(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1041), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1042), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1108), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT122), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1348), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1059), .A2(G2067), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n619), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1114), .A2(KEYINPUT122), .A3(new_n1118), .A4(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1113), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1114), .A2(KEYINPUT61), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(new_n1070), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1113), .B1(new_n1123), .B2(new_n1114), .ZN(new_n1124));
  INV_X1    g699(.A(G1996), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1009), .A2(new_n1125), .A3(new_n1013), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  AOI22_X1  g703(.A1(new_n1126), .A2(new_n1127), .B1(new_n1059), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1041), .A2(KEYINPUT121), .A3(new_n1125), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n559), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT59), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1116), .A2(new_n619), .A3(new_n1117), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n619), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1124), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1072), .A2(G301), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1078), .A2(KEYINPUT54), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT54), .B1(new_n1078), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1122), .A2(new_n1139), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1082), .A2(new_n1103), .A3(new_n1104), .A4(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1017), .A2(new_n1000), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n773), .B(G1996), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n797), .B(G2067), .Z(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n753), .ZN(new_n1151));
  INV_X1    g726(.A(new_n755), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1147), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1146), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1147), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n797), .A2(G2067), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT48), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1160), .A2(G1986), .A3(G290), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1156), .A2(new_n1147), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1165), .A2(new_n1164), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1160), .B1(new_n773), .B2(new_n1149), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT126), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1147), .A2(new_n1125), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT46), .Z(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT127), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT47), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1168), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1175), .B2(new_n1174), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(new_n993), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n684), .A2(G319), .A3(new_n665), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G229), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n910), .A3(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


