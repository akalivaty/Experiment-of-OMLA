//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1179, new_n1180, new_n1181, new_n1182, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G50), .A2(G226), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT66), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n215), .A2(new_n216), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G97), .A2(G257), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n211), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT69), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n232), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT70), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n255), .A3(new_n252), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G226), .A3(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n251), .B(G274), .C1(G41), .C2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G222), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G223), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n250), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n265), .B(new_n266), .C1(G77), .C2(new_n261), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT71), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n257), .A2(new_n268), .A3(new_n258), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n225), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n251), .B2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n202), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n226), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(G20), .B2(new_n203), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n273), .A2(new_n225), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n276), .B(new_n279), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n272), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n270), .A2(G179), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n288), .B(KEYINPUT9), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT73), .B(G200), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n270), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n260), .A2(G190), .A3(new_n267), .A4(new_n269), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n292), .A2(new_n298), .A3(new_n294), .A4(new_n295), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n291), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  OAI211_X1 g0102(.A(G226), .B(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(G232), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n266), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n254), .A2(G238), .A3(new_n256), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n258), .B(KEYINPUT74), .Z(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(G179), .A3(new_n313), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n318), .A3(G169), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n284), .A2(new_n202), .B1(new_n226), .B2(G68), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n281), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n274), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT11), .ZN(new_n325));
  INV_X1    g0125(.A(G13), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G1), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G20), .A3(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT12), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT12), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(G68), .B2(new_n275), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n314), .B2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n311), .A2(G190), .A3(new_n313), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n261), .A2(G232), .A3(new_n263), .ZN(new_n342));
  INV_X1    g0142(.A(G107), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n261), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n266), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n254), .A2(G244), .A3(new_n256), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n258), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n271), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n347), .A2(G179), .ZN(new_n349));
  INV_X1    g0149(.A(new_n280), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT15), .B(G87), .Z(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n281), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n274), .B1(new_n322), .B2(new_n278), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n275), .A2(G77), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT72), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT72), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n348), .B(new_n349), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n300), .A2(new_n334), .A3(new_n340), .A4(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n301), .A2(new_n302), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n362), .B2(new_n226), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n301), .A2(new_n302), .A3(new_n364), .A4(G20), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n283), .A2(G159), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n328), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n201), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n367), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n364), .B1(new_n261), .B2(G20), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n362), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n328), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(new_n367), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n377), .A3(new_n274), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n350), .A2(new_n277), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n350), .B2(new_n275), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  OAI211_X1 g0182(.A(G223), .B(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n261), .A2(new_n385), .A3(G223), .A4(new_n263), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n261), .A2(G226), .A3(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n384), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n266), .ZN(new_n390));
  INV_X1    g0190(.A(G232), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n258), .B1(new_n253), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n382), .B1(new_n394), .B2(G179), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n271), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n389), .B2(new_n266), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(KEYINPUT77), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n381), .A2(new_n395), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n399), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT77), .B1(new_n397), .B2(new_n398), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(KEYINPUT18), .A3(new_n381), .A4(new_n396), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n397), .A2(G200), .ZN(new_n408));
  AOI211_X1 g0208(.A(G190), .B(new_n392), .C1(new_n389), .C2(new_n266), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n378), .B(new_n380), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n397), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G200), .B2(new_n397), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n378), .A4(new_n380), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n359), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n347), .A2(new_n413), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n347), .A2(new_n293), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n357), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n361), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(G264), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n426));
  OAI211_X1 g0226(.A(G257), .B(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n427));
  OR2_X1    g0227(.A1(KEYINPUT3), .A2(G33), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT3), .A2(G33), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(G303), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n266), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1), .ZN(new_n434));
  INV_X1    g0234(.A(G41), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G41), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G274), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(G270), .A3(new_n250), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n432), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n327), .A2(G20), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n251), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n287), .A2(G116), .A3(new_n277), .A4(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n273), .A2(new_n225), .B1(G20), .B2(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n226), .C1(G33), .C2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT20), .B1(new_n449), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n446), .B(new_n448), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n444), .A2(G169), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT21), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n444), .A2(G200), .ZN(new_n459));
  INV_X1    g0259(.A(new_n455), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n432), .A2(G190), .A3(new_n442), .A4(new_n443), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n439), .A2(new_n250), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n266), .A2(new_n431), .B1(new_n463), .B2(G270), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n455), .A3(G179), .A4(new_n442), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n444), .A2(KEYINPUT21), .A3(new_n455), .A4(G169), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n458), .A2(new_n462), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n226), .B(G87), .C1(new_n301), .C2(new_n302), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT22), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(KEYINPUT82), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n261), .A2(new_n226), .A3(G87), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n226), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n226), .B2(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n343), .A2(KEYINPUT23), .A3(G20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n471), .A2(new_n474), .A3(new_n477), .A4(new_n481), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT83), .B(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n469), .A2(new_n470), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  INV_X1    g0285(.A(new_n483), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n474), .A3(new_n477), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n274), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G257), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n489));
  OAI211_X1 g0289(.A(G250), .B(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G294), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n266), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n439), .A2(G264), .A3(new_n250), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n442), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n287), .A2(new_n277), .A3(new_n447), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n327), .A2(G20), .A3(new_n343), .ZN(new_n500));
  XOR2_X1   g0300(.A(new_n500), .B(KEYINPUT25), .Z(new_n501));
  NAND4_X1  g0301(.A1(new_n488), .A2(new_n496), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n495), .A2(new_n413), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n352), .A2(new_n277), .ZN(new_n505));
  INV_X1    g0305(.A(G87), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n281), .B2(new_n451), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n261), .A2(new_n226), .A3(G68), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n508), .C1(new_n281), .C2(new_n451), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n226), .B1(new_n305), .B2(new_n508), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n511), .A3(new_n513), .A4(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n505), .B(new_n507), .C1(new_n518), .C2(new_n274), .ZN(new_n519));
  OR2_X1    g0319(.A1(G238), .A2(G1698), .ZN(new_n520));
  OAI221_X1 g0320(.A(new_n520), .B1(G244), .B2(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n250), .B1(new_n521), .B2(new_n475), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n434), .A2(G274), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n433), .B2(G1), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n251), .A2(KEYINPUT80), .A3(G45), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n250), .A2(new_n526), .A3(G250), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n522), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  INV_X1    g0331(.A(G244), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n428), .A2(new_n429), .B1(new_n532), .B2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n476), .B1(new_n533), .B2(new_n520), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n523), .B(new_n528), .C1(new_n534), .C2(new_n250), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n293), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n519), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n398), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n505), .B1(new_n518), .B2(new_n274), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n498), .A2(new_n352), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n271), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n488), .A2(new_n499), .A3(new_n501), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n495), .A2(new_n271), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n266), .A2(new_n492), .B1(new_n463), .B2(G264), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n398), .A3(new_n442), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n468), .A2(new_n504), .A3(new_n544), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT79), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT6), .ZN(new_n553));
  AND2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n515), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n343), .A2(KEYINPUT6), .A3(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n226), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n284), .A2(new_n322), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n558), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n343), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n553), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT78), .B(new_n560), .C1(new_n563), .C2(new_n226), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n363), .B2(new_n365), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n274), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n278), .A2(new_n451), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n498), .A2(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(new_n263), .C1(new_n301), .C2(new_n302), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n450), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n266), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n441), .B1(new_n463), .B2(G257), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n271), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n398), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n570), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n566), .A2(new_n274), .B1(new_n451), .B2(new_n278), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(G200), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(G190), .A3(new_n578), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n569), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n551), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n583), .A2(new_n551), .A3(new_n587), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n550), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n425), .A2(new_n591), .ZN(G372));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  INV_X1    g0393(.A(new_n333), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n318), .B1(new_n314), .B2(G169), .ZN(new_n595));
  AOI211_X1 g0395(.A(KEYINPUT14), .B(new_n271), .C1(new_n311), .C2(new_n313), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n597), .B2(new_n317), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n314), .A2(G200), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n594), .A3(new_n337), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n360), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n593), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n334), .B(KEYINPUT85), .C1(new_n601), .C2(new_n360), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n418), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n407), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n297), .A2(new_n299), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n291), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n543), .B(new_n537), .C1(new_n502), .C2(new_n503), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n583), .A2(new_n587), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n549), .A2(KEYINPUT84), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n545), .A2(new_n613), .A3(new_n546), .A4(new_n548), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n458), .A2(new_n465), .A3(new_n466), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n610), .B(new_n611), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n543), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n584), .A2(new_n569), .B1(new_n271), .B2(new_n579), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n544), .A2(KEYINPUT26), .A3(new_n619), .A4(new_n582), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n537), .A2(new_n543), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n583), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n425), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n608), .A2(new_n626), .ZN(G369));
  NOR3_X1   g0427(.A1(new_n326), .A2(G1), .A3(G20), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT27), .ZN(new_n629));
  OR3_X1    g0429(.A1(new_n628), .A2(KEYINPUT86), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G213), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n628), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT86), .B1(new_n628), .B2(new_n629), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G343), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n460), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n467), .B2(new_n638), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n545), .A2(new_n636), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n504), .A2(new_n549), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n616), .A2(new_n637), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n643), .B(new_n644), .C1(new_n549), .C2(new_n637), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n502), .A2(new_n503), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n615), .B2(new_n637), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(G399));
  NOR2_X1   g0451(.A1(new_n516), .A2(G116), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n209), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n653), .A2(new_n655), .A3(new_n251), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  INV_X1    g0459(.A(new_n655), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n658), .B(new_n659), .C1(new_n228), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT28), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT89), .B1(new_n647), .B2(new_n616), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n458), .A2(new_n466), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n549), .A3(new_n665), .A4(new_n465), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n663), .A2(new_n611), .A3(new_n610), .A4(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n636), .B1(new_n624), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT29), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI211_X1 g0470(.A(KEYINPUT29), .B(new_n636), .C1(new_n617), .C2(new_n624), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n609), .A2(new_n647), .A3(new_n467), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n583), .A2(new_n551), .A3(new_n587), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n673), .B(new_n637), .C1(new_n588), .C2(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n444), .A2(new_n535), .A3(new_n398), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT30), .A3(new_n581), .A4(new_n547), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n530), .A2(G179), .A3(new_n442), .A4(new_n464), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n577), .A2(new_n547), .A3(new_n578), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(G179), .B1(new_n547), .B2(new_n442), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n535), .A3(new_n444), .A4(new_n579), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n636), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n636), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n675), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n672), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n662), .B1(new_n693), .B2(G1), .ZN(G364));
  XOR2_X1   g0494(.A(new_n641), .B(KEYINPUT90), .Z(new_n695));
  NOR2_X1   g0495(.A1(new_n326), .A2(G20), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n251), .B1(new_n696), .B2(G45), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n655), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n695), .B(new_n700), .C1(G330), .C2(new_n640), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n654), .A2(new_n362), .ZN(new_n702));
  NAND2_X1  g0502(.A1(G355), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n654), .A2(new_n261), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n247), .B2(new_n433), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n228), .A2(G45), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n703), .B1(G116), .B2(new_n209), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G13), .A2(G33), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n225), .B1(G20), .B2(new_n271), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n226), .A2(G190), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G179), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G159), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT32), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n362), .B1(new_n718), .B2(KEYINPUT32), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n226), .A2(new_n413), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n293), .A2(new_n398), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G87), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n293), .A2(new_n398), .A3(new_n714), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G107), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n719), .A2(new_n720), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n398), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n714), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(G58), .A2(new_n731), .B1(new_n733), .B2(G77), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n226), .B1(new_n715), .B2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n226), .A2(new_n398), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n734), .B1(new_n451), .B2(new_n735), .C1(new_n328), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n737), .A2(new_n413), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n728), .B(new_n740), .C1(G50), .C2(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G283), .A2(new_n726), .B1(new_n723), .B2(G303), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n743), .B(new_n362), .C1(new_n744), .C2(new_n730), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n738), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  INV_X1    g0551(.A(new_n741), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(new_n750), .B2(new_n732), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n717), .A2(G329), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n745), .A2(new_n753), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n711), .B1(new_n742), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n710), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n713), .B(new_n758), .C1(new_n640), .C2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n701), .B1(new_n700), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT91), .ZN(G396));
  NAND2_X1  g0562(.A1(new_n625), .A2(new_n637), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n360), .A2(new_n636), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n636), .B1(new_n358), .B2(new_n359), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n423), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n360), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n764), .B1(new_n767), .B2(new_n360), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n625), .A2(new_n637), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G330), .A3(new_n690), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(new_n691), .A3(new_n772), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n700), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n739), .A2(new_n777), .B1(new_n735), .B2(new_n451), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n261), .B(new_n778), .C1(G303), .C2(new_n741), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n723), .A2(G107), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G294), .A2(new_n731), .B1(new_n733), .B2(G116), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n725), .A2(new_n506), .B1(new_n750), .B2(new_n716), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G137), .A2(new_n741), .B1(new_n738), .B2(G150), .ZN(new_n785));
  INV_X1    g0585(.A(G143), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n785), .B1(new_n786), .B2(new_n730), .C1(new_n787), .C2(new_n732), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT93), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT34), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n261), .B1(new_n791), .B2(new_n716), .C1(new_n722), .C2(new_n202), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n790), .B(new_n793), .C1(new_n328), .C2(new_n725), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n735), .A2(new_n368), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n784), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n711), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n711), .A2(new_n708), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(G77), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n771), .A2(new_n709), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n699), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n776), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G384));
  INV_X1    g0607(.A(KEYINPUT38), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT96), .ZN(new_n809));
  INV_X1    g0609(.A(new_n400), .ZN(new_n810));
  INV_X1    g0610(.A(new_n634), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n381), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n410), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n809), .B(KEYINPUT37), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n417), .B1(new_n402), .B2(new_n406), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n812), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT37), .B1(new_n810), .B2(new_n813), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT37), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n400), .A2(new_n818), .A3(new_n410), .A4(new_n812), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n817), .A2(KEYINPUT96), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n808), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n812), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n419), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n817), .A2(KEYINPUT96), .A3(new_n819), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n823), .A2(KEYINPUT38), .A3(new_n824), .A4(new_n814), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n821), .A2(KEYINPUT39), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n817), .A2(new_n819), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n812), .B1(new_n407), .B2(new_n418), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n334), .A2(new_n636), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n407), .A2(new_n811), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n333), .A2(new_n636), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n340), .B2(new_n334), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n600), .A2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n598), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n764), .B(KEYINPUT95), .Z(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n772), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n821), .A2(new_n825), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n835), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n425), .B1(new_n670), .B2(new_n671), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n608), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n846), .B(new_n848), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n600), .A2(KEYINPUT75), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n333), .B(new_n636), .C1(new_n852), .C2(new_n320), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n334), .A2(new_n600), .A3(new_n837), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n636), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n688), .B1(new_n684), .B2(new_n636), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n675), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n859), .A3(new_n771), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n825), .B2(new_n821), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT98), .B1(new_n861), .B2(KEYINPUT40), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n855), .A2(new_n859), .A3(new_n771), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n844), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT98), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n769), .B1(new_n853), .B2(new_n854), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n859), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n831), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n825), .A2(new_n830), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n863), .A2(new_n872), .A3(KEYINPUT99), .A4(KEYINPUT40), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n862), .A2(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n425), .A3(new_n859), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n873), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT98), .B(KEYINPUT40), .C1(new_n844), .C2(new_n863), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n876), .B(G330), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G330), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n675), .B2(new_n858), .ZN(new_n881));
  AND4_X1   g0681(.A1(new_n300), .A2(new_n334), .A3(new_n340), .A4(new_n360), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n419), .A2(new_n424), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n849), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n251), .B2(new_n696), .ZN(new_n888));
  INV_X1    g0688(.A(new_n563), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n445), .B1(new_n889), .B2(KEYINPUT35), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n227), .C1(KEYINPUT35), .C2(new_n889), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  OAI21_X1  g0692(.A(G77), .B1(new_n368), .B2(new_n328), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n893), .A2(new_n228), .B1(G50), .B2(new_n328), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n326), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n892), .A3(new_n895), .ZN(G367));
  INV_X1    g0696(.A(new_n704), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n712), .B1(new_n209), .B2(new_n353), .C1(new_n240), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n726), .A2(G77), .ZN(new_n899));
  AOI22_X1  g0699(.A1(G150), .A2(new_n731), .B1(new_n717), .B2(G137), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n901), .B1(new_n202), .B2(new_n732), .C1(new_n786), .C2(new_n752), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n722), .A2(new_n368), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n739), .A2(new_n787), .B1(new_n735), .B2(new_n328), .ZN(new_n904));
  NOR4_X1   g0704(.A1(new_n902), .A2(new_n362), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n723), .A2(KEYINPUT46), .A3(G116), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT104), .Z(new_n907));
  AOI211_X1 g0707(.A(new_n261), .B(new_n907), .C1(G97), .C2(new_n726), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n732), .A2(new_n777), .B1(new_n735), .B2(new_n343), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n908), .B1(KEYINPUT103), .B2(new_n909), .C1(new_n754), .C2(new_n739), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT46), .B1(new_n723), .B2(G116), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT105), .Z(new_n912));
  AOI22_X1  g0712(.A1(new_n909), .A2(KEYINPUT103), .B1(G303), .B2(new_n731), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n746), .B2(new_n716), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n741), .A2(G311), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n905), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT47), .ZN(new_n918));
  INV_X1    g0718(.A(new_n711), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n699), .B(new_n898), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n519), .A2(new_n637), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n543), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n544), .B2(new_n921), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT100), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n924), .A2(new_n710), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n570), .A2(new_n636), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n611), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n619), .A2(new_n582), .A3(new_n636), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n649), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT42), .Z(new_n932));
  OAI21_X1  g0732(.A(new_n583), .B1(new_n928), .B2(new_n549), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n637), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT43), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n924), .A2(new_n936), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT101), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n940), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n646), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n930), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n942), .A2(new_n945), .A3(new_n930), .A4(new_n943), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n655), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n649), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n645), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n695), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n646), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n692), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT102), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n650), .A2(new_n956), .A3(new_n930), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n956), .B1(new_n650), .B2(new_n930), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n650), .A2(new_n930), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT44), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n950), .B1(new_n965), .B2(new_n692), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n697), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n926), .B1(new_n949), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(G387));
  OAI221_X1 g0769(.A(new_n362), .B1(new_n751), .B2(new_n716), .C1(new_n725), .C2(new_n445), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G311), .A2(new_n738), .B1(new_n741), .B2(G322), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT107), .Z(new_n972));
  INV_X1    g0772(.A(G303), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n973), .B2(new_n732), .C1(new_n746), .C2(new_n730), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n777), .B2(new_n735), .C1(new_n754), .C2(new_n722), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT49), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT49), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n732), .A2(new_n328), .B1(new_n716), .B2(new_n282), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n722), .A2(new_n322), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G159), .C2(new_n741), .ZN(new_n982));
  INV_X1    g0782(.A(new_n735), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n352), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n202), .B2(new_n730), .C1(new_n280), .C2(new_n739), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n362), .B(new_n986), .C1(G97), .C2(new_n726), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n711), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n643), .B(new_n710), .C1(new_n549), .C2(new_n637), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n653), .A2(new_n702), .B1(new_n343), .B2(new_n654), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n237), .A2(G45), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n280), .A2(KEYINPUT50), .A3(G50), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT50), .B1(new_n280), .B2(G50), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n992), .A2(new_n993), .A3(new_n433), .A4(new_n652), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n328), .A2(new_n322), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n704), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT106), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n712), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n988), .A2(new_n699), .A3(new_n989), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n954), .A2(new_n692), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n655), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1000), .B1(new_n697), .B2(new_n954), .C1(new_n955), .C2(new_n1002), .ZN(G393));
  NAND2_X1  g0803(.A1(new_n964), .A2(new_n945), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n960), .A2(new_n962), .A3(new_n646), .A4(new_n963), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n955), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1006), .A2(new_n965), .A3(new_n660), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT108), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n698), .A3(new_n1005), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n741), .A2(G317), .B1(new_n731), .B2(G311), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT52), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G322), .B2(new_n717), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n733), .A2(G294), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n261), .B1(new_n723), .B2(G283), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n738), .A2(G303), .B1(G116), .B2(new_n983), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1015), .A2(new_n727), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n741), .A2(G150), .B1(new_n731), .B2(G159), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT51), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G87), .B2(new_n726), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n362), .B1(new_n723), .B2(G68), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G77), .B2(new_n983), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n786), .B2(new_n716), .C1(new_n280), .C2(new_n732), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n739), .A2(new_n202), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1017), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n711), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n712), .B1(new_n451), .B2(new_n209), .C1(new_n244), .C2(new_n897), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n928), .A2(new_n710), .A3(new_n929), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n699), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1007), .A2(new_n1008), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1008), .B1(new_n1007), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(G390));
  INV_X1    g0834(.A(new_n843), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT110), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n834), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT110), .B1(new_n843), .B2(new_n833), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n832), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n833), .B(KEYINPUT109), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n668), .A2(new_n771), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(new_n842), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n872), .B(new_n1040), .C1(new_n1042), .C2(new_n841), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n855), .A2(new_n859), .A3(G330), .A4(new_n771), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT111), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT111), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n869), .A2(new_n1047), .A3(G330), .A4(new_n859), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  AND4_X1   g0850(.A1(G330), .A2(new_n690), .A3(new_n855), .A4(new_n771), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1039), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n690), .A2(G330), .A3(new_n771), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n841), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1046), .A2(new_n1055), .A3(new_n1048), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n772), .A2(new_n842), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n690), .A2(new_n855), .A3(G330), .A4(new_n771), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n881), .A2(new_n771), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1042), .B(new_n1059), .C1(new_n1060), .C2(new_n855), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n884), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n425), .A2(KEYINPUT112), .A3(new_n881), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n608), .A2(new_n847), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1053), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1068), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n660), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n832), .A2(new_n708), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n350), .B2(new_n799), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n261), .B1(new_n725), .B2(new_n202), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n717), .A2(G125), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n983), .A2(G159), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n738), .A2(G137), .B1(new_n731), .B2(G132), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n722), .A2(new_n282), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT53), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT54), .B(G143), .Z(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT113), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1088), .A2(new_n733), .B1(G128), .B2(new_n741), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n724), .B1(new_n445), .B2(new_n730), .C1(new_n777), .C2(new_n752), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G294), .B2(new_n717), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n738), .A2(G107), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n726), .A2(G68), .B1(G77), .B2(new_n983), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n261), .B1(new_n733), .B2(G97), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n919), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1075), .A2(new_n700), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1053), .B2(new_n697), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1073), .A2(new_n1101), .ZN(G378));
  OAI22_X1  g0902(.A1(new_n739), .A2(new_n791), .B1(new_n735), .B2(new_n282), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G125), .B2(new_n741), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n733), .A2(G137), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1088), .A2(new_n723), .B1(G128), .B2(new_n731), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n435), .ZN(new_n1109));
  AOI211_X1 g0909(.A(G33), .B(new_n1109), .C1(G124), .C2(new_n717), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(KEYINPUT59), .B2(new_n1107), .C1(new_n787), .C2(new_n725), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n202), .B1(new_n301), .B2(G41), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n981), .B1(G97), .B2(new_n738), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n726), .A2(G58), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n777), .C2(new_n716), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n735), .A2(new_n328), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n752), .A2(new_n445), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n362), .B1(new_n353), .B2(new_n732), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n435), .C1(new_n343), .C2(new_n730), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT58), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1111), .A2(new_n1112), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n288), .A2(new_n811), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n300), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n300), .A2(new_n1123), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1129), .A2(KEYINPUT116), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT116), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n699), .B1(new_n919), .B2(new_n1122), .C1(new_n1134), .C2(new_n709), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n202), .B2(new_n798), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT117), .B1(new_n879), .B2(new_n1133), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n874), .A2(new_n1134), .A3(new_n1138), .A4(G330), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n879), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n846), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n846), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1137), .A2(new_n1140), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1136), .B1(new_n1145), .B2(new_n698), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n655), .B1(new_n1148), .B2(KEYINPUT57), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT57), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1150), .B(new_n1147), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1146), .B1(new_n1149), .B2(new_n1151), .ZN(G375));
  OAI21_X1  g0952(.A(new_n699), .B1(new_n799), .B2(G68), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(KEYINPUT118), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n261), .B1(new_n282), .B2(new_n732), .C1(new_n722), .C2(new_n787), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1088), .A2(new_n738), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n983), .A2(G50), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G137), .A2(new_n731), .B1(new_n717), .B2(G128), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1156), .A2(new_n1114), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1155), .B(new_n1159), .C1(G132), .C2(new_n741), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G283), .A2(new_n731), .B1(new_n733), .B2(G107), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n899), .C1(new_n973), .C2(new_n716), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n261), .B1(new_n738), .B2(G116), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1163), .B(new_n984), .C1(new_n754), .C2(new_n752), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G97), .C2(new_n723), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n711), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1153), .A2(KEYINPUT118), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1154), .B(new_n1168), .C1(new_n841), .C2(new_n708), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1062), .B2(new_n698), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1058), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n950), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1071), .B2(new_n1172), .ZN(G381));
  XOR2_X1   g0973(.A(G375), .B(KEYINPUT119), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(G378), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n968), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1176), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n806), .A3(new_n1177), .ZN(G407));
  NAND2_X1  g0978(.A1(new_n635), .A2(G213), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT120), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n631), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(G407), .ZN(G409));
  XNOR2_X1  g0983(.A(G393), .B(G396), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1176), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n968), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(G390), .A2(G387), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1176), .A3(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1187), .A2(KEYINPUT126), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT126), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT61), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT124), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n655), .A3(new_n1068), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1058), .A2(KEYINPUT60), .A3(new_n1061), .A4(new_n1066), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n855), .B1(new_n881), .B2(new_n771), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1051), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1057), .A2(new_n1056), .B1(new_n1202), .B2(new_n1042), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1203), .A2(new_n1204), .A3(KEYINPUT60), .A4(new_n1066), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1200), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1170), .B1(new_n1198), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(G384), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n660), .B1(new_n1171), .B2(new_n1196), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1209), .A2(new_n1200), .A3(new_n1068), .A4(new_n1205), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n806), .A3(new_n1170), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(G2897), .A3(new_n1181), .A4(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT123), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n635), .A2(G213), .A3(G2897), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1210), .A2(new_n806), .A3(new_n1170), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n806), .B1(new_n1210), .B2(new_n1170), .ZN(new_n1218));
  OAI211_X1 g1018(.A(KEYINPUT122), .B(new_n1215), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1195), .B1(new_n1213), .B2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1223), .A2(KEYINPUT123), .A3(G2897), .A4(new_n1181), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1212), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1219), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1231), .A3(KEYINPUT124), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1222), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1146), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1148), .A2(new_n950), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1146), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1073), .A2(new_n1101), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1181), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1194), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1179), .A3(new_n1214), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1223), .A2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1242), .A2(new_n1243), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1193), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1227), .A2(new_n1231), .A3(KEYINPUT124), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT124), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1222), .A2(KEYINPUT125), .A3(new_n1232), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1241), .A2(new_n1179), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1223), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1242), .A2(new_n1254), .B1(new_n1190), .B2(new_n1187), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1246), .A2(new_n1258), .ZN(G405));
  AND2_X1   g1059(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1150), .B1(new_n1260), .B2(new_n1147), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1148), .A2(KEYINPUT57), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n655), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G378), .B1(new_n1263), .B2(new_n1146), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1234), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1214), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G375), .A2(new_n1237), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1223), .A3(new_n1234), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1193), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1193), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1266), .A2(new_n1193), .A3(KEYINPUT127), .A4(new_n1268), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1271), .A2(new_n1274), .A3(new_n1275), .ZN(G402));
endmodule


