//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n203), .A2(G50), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT66), .Z(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n210), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT67), .Z(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G50), .B2(G226), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n215), .B(new_n230), .C1(new_n211), .C2(new_n214), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT13), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G226), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(G1698), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(G33), .B2(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n251), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n264), .A2(G238), .A3(new_n249), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n247), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n256), .B2(new_n257), .ZN(new_n268));
  NOR4_X1   g0068(.A1(new_n268), .A2(KEYINPUT13), .A3(new_n265), .A4(new_n251), .ZN(new_n269));
  OAI21_X1  g0069(.A(G169), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT14), .ZN(new_n271));
  INV_X1    g0071(.A(new_n251), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n254), .A2(new_n255), .B1(G33), .B2(G97), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n266), .B(new_n272), .C1(new_n264), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n258), .A2(new_n260), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n276), .A2(new_n247), .A3(new_n272), .A4(new_n266), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G179), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n277), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT14), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(G169), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n271), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n262), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(G77), .B1(new_n284), .B2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(G20), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G68), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n259), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n248), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G68), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G68), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT11), .B1(new_n287), .B2(new_n289), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n275), .A2(G190), .A3(new_n277), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n275), .B2(new_n277), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT72), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n279), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n301), .A3(new_n307), .A4(new_n298), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(G222), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G223), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n260), .C1(G77), .C2(new_n255), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n264), .A2(new_n249), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n272), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(G179), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT8), .B(G58), .Z(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n283), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  INV_X1    g0130(.A(new_n284), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G50), .ZN(new_n333));
  INV_X1    g0133(.A(new_n294), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n332), .A2(new_n289), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n291), .A2(G50), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n326), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n310), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT15), .A2(G87), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT15), .A2(G87), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT15), .A2(G87), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT69), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n349), .A3(new_n283), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT70), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G20), .A2(G77), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT70), .A4(new_n283), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n327), .A2(new_n284), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n289), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n334), .A2(new_n226), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n291), .A2(G77), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G238), .A2(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n255), .B(new_n361), .C1(new_n253), .C2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n260), .C1(G107), .C2(new_n255), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n320), .A2(G244), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n272), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G169), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n363), .A2(G179), .A3(new_n272), .A4(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n356), .A2(new_n289), .B1(new_n226), .B2(new_n334), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT71), .B(G200), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n363), .A2(G190), .A3(new_n272), .A4(new_n364), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n370), .A2(new_n372), .A3(new_n359), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n342), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n337), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT9), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n325), .A2(new_n371), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n325), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT9), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n337), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n380), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n382), .A2(new_n377), .A3(new_n384), .A4(new_n378), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n327), .A2(new_n294), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n327), .B2(new_n291), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT73), .B1(new_n311), .B2(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n312), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n311), .A2(KEYINPUT73), .A3(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n321), .A2(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n317), .A2(new_n315), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n260), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n320), .A2(G232), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n399), .A2(new_n381), .A3(new_n400), .A4(new_n272), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n264), .B1(new_n396), .B2(new_n397), .ZN(new_n402));
  INV_X1    g0202(.A(new_n400), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n402), .A2(new_n403), .A3(new_n251), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n401), .B1(new_n404), .B2(G200), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n255), .B2(G20), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n311), .A2(G33), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT7), .B(new_n286), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT74), .B1(new_n411), .B2(G68), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  INV_X1    g0213(.A(G68), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n407), .C2(new_n410), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G58), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n414), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(new_n202), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(G20), .B1(G159), .B2(new_n284), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT16), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n422));
  OAI21_X1  g0222(.A(G68), .B1(new_n422), .B2(new_n406), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(KEYINPUT3), .B2(new_n262), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n393), .B1(new_n425), .B2(new_n408), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n286), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n428));
  OAI211_X1 g0228(.A(KEYINPUT16), .B(new_n420), .C1(new_n423), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n289), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n390), .B(new_n405), .C1(new_n421), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n289), .ZN(new_n434));
  INV_X1    g0234(.A(new_n420), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n414), .B1(new_n427), .B2(KEYINPUT7), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n422), .A2(new_n406), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n255), .A2(new_n406), .A3(G20), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT7), .B1(new_n314), .B2(new_n286), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n413), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n411), .A2(KEYINPUT74), .A3(G68), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n420), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(KEYINPUT17), .A3(new_n390), .A4(new_n405), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n433), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(new_n390), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n439), .B2(new_n447), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n404), .A2(new_n338), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n402), .A2(new_n403), .A3(new_n455), .A4(new_n251), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n451), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n390), .B1(new_n421), .B2(new_n430), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n404), .A2(G179), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n338), .B2(new_n404), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(KEYINPUT18), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n388), .A2(new_n450), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n375), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n248), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n294), .A2(new_n466), .A3(new_n259), .A4(new_n288), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n334), .A2(KEYINPUT25), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT25), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n294), .B2(G107), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n468), .A2(G107), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n218), .A2(G20), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n312), .A3(new_n313), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT23), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n286), .B2(G107), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n475), .A2(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n392), .A2(KEYINPUT22), .A3(new_n474), .A4(new_n393), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n283), .A2(G116), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT24), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n480), .A2(new_n481), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT79), .B1(new_n487), .B2(new_n289), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n434), .C1(new_n484), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n473), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G1), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G264), .A3(new_n264), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n248), .A2(G45), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n263), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n494), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G274), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n221), .A2(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n219), .A2(new_n315), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n392), .A2(new_n393), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G294), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n504), .B1(new_n260), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G169), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n455), .B2(new_n510), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n491), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n260), .ZN(new_n514));
  INV_X1    g0314(.A(new_n504), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT80), .B1(new_n516), .B2(G190), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n303), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n519), .A3(new_n381), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n473), .C1(new_n488), .C2(new_n490), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n294), .B2(G97), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n294), .A2(new_n524), .A3(G97), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n525), .A2(new_n527), .B1(new_n468), .B2(G97), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT75), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n411), .B2(G107), .ZN(new_n530));
  AOI211_X1 g0330(.A(KEYINPUT75), .B(new_n469), .C1(new_n407), .C2(new_n410), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n532), .A2(new_n220), .A3(G107), .ZN(new_n533));
  XNOR2_X1  g0333(.A(G97), .B(G107), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n535), .A2(new_n286), .B1(new_n226), .B2(new_n331), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n528), .B1(new_n537), .B2(new_n434), .ZN(new_n538));
  INV_X1    g0338(.A(new_n393), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n312), .B2(new_n391), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT4), .B1(new_n540), .B2(G244), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n315), .A2(KEYINPUT4), .A3(G244), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n543), .B1(new_n255), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n255), .B2(G250), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n315), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n260), .B1(new_n541), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n502), .A2(new_n260), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n503), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n338), .ZN(new_n554));
  INV_X1    g0354(.A(new_n552), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n312), .A2(new_n313), .A3(G250), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n315), .B1(new_n556), .B2(KEYINPUT4), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n542), .B1(new_n314), .B2(new_n544), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n547), .B1(new_n426), .B2(new_n227), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n555), .B1(new_n561), .B2(new_n260), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n455), .A3(new_n503), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n538), .A2(new_n554), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n528), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n411), .A2(G107), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g0367(.A(new_n536), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n411), .A2(new_n529), .A3(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n565), .B1(new_n570), .B2(new_n289), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n562), .A2(G190), .A3(new_n503), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n553), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT19), .B1(new_n283), .B2(G97), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n218), .A2(new_n220), .A3(new_n469), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n257), .A2(new_n286), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n578), .B2(KEYINPUT19), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n392), .A2(new_n286), .A3(G68), .A4(new_n393), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n434), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n347), .A2(new_n349), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n294), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n467), .A2(new_n218), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G116), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n227), .A2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G238), .B2(G1698), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n426), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G238), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n227), .B2(G1698), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n392), .A2(new_n593), .A3(new_n393), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(KEYINPUT77), .A3(new_n586), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n260), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n260), .A2(new_n493), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(G250), .B1(G274), .B2(new_n493), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n596), .A2(new_n381), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n371), .B1(new_n596), .B2(new_n598), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n585), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n594), .A2(KEYINPUT77), .A3(new_n586), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT77), .B1(new_n594), .B2(new_n586), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n603), .A3(new_n264), .ZN(new_n604));
  INV_X1    g0404(.A(new_n598), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n338), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n596), .A2(new_n455), .A3(new_n598), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n581), .A2(new_n583), .ZN(new_n608));
  INV_X1    g0408(.A(new_n582), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n467), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n564), .A2(new_n574), .A3(new_n601), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G264), .A2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n221), .B2(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n392), .A2(new_n393), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n314), .A2(G303), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n260), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n497), .A2(G270), .A3(new_n264), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n503), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n338), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n542), .B(new_n286), .C1(G33), .C2(new_n220), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G20), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n289), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n623), .A2(KEYINPUT20), .A3(new_n289), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT78), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n294), .A2(G116), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n468), .B2(G116), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n630), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n622), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n622), .B(KEYINPUT21), .C1(new_n634), .C2(new_n635), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(new_n633), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT78), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n264), .B1(new_n615), .B2(new_n616), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n644), .A2(new_n620), .A3(new_n455), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n618), .A2(new_n621), .A3(G190), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n644), .B2(new_n620), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n641), .A2(new_n647), .A3(new_n642), .A4(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n638), .A2(new_n639), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n523), .A2(new_n612), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n465), .A2(new_n651), .ZN(G372));
  NAND3_X1  g0452(.A1(new_n638), .A2(new_n639), .A3(new_n646), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n491), .B2(new_n512), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n564), .B(new_n574), .C1(new_n491), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n585), .A2(KEYINPUT81), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT81), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n581), .A2(new_n583), .A3(new_n658), .A4(new_n584), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n657), .A2(new_n659), .B1(new_n599), .B2(new_n600), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n611), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n654), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n601), .A2(new_n611), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n663), .B2(new_n564), .ZN(new_n664));
  AOI21_X1  g0464(.A(G169), .B1(new_n562), .B2(new_n503), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n455), .A2(new_n550), .A3(new_n503), .A4(new_n552), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n571), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n611), .A4(new_n660), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(new_n669), .A3(new_n611), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n465), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n387), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT82), .B1(new_n385), .B2(new_n387), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n369), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n309), .A2(new_n675), .B1(new_n299), .B2(new_n282), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n433), .A2(new_n449), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n463), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n341), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(G369));
  AND4_X1   g0480(.A1(new_n638), .A2(new_n649), .A3(new_n639), .A4(new_n646), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT84), .ZN(new_n682));
  INV_X1    g0482(.A(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G20), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n248), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT83), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT83), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n685), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(G213), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n643), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n682), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n653), .B2(new_n695), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n513), .A2(new_n522), .ZN(new_n700));
  INV_X1    g0500(.A(new_n491), .ZN(new_n701));
  INV_X1    g0501(.A(new_n694), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n513), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n694), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n653), .A2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n709), .C1(new_n513), .C2(new_n694), .ZN(G399));
  NOR2_X1   g0510(.A1(new_n576), .A2(G116), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT85), .Z(new_n712));
  INV_X1    g0512(.A(new_n213), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(G1), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n209), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n702), .B1(new_n662), .B2(new_n670), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT88), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(KEYINPUT88), .B(new_n702), .C1(new_n662), .C2(new_n670), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT29), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(new_n611), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n667), .A2(new_n611), .A3(new_n660), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n667), .A2(new_n668), .A3(new_n601), .A4(new_n611), .ZN(new_n729));
  INV_X1    g0529(.A(new_n661), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n704), .B2(new_n653), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n656), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n725), .B1(new_n732), .B2(new_n702), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n724), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT87), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n596), .A2(new_n598), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n455), .B1(new_n644), .B2(new_n620), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n553), .A2(new_n736), .A3(new_n516), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT86), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n562), .A2(new_n645), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n596), .A2(new_n510), .A3(new_n598), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n645), .A2(new_n550), .A3(new_n552), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n604), .A2(new_n605), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT30), .A4(new_n510), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n737), .B1(new_n596), .B2(new_n598), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT86), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n516), .A4(new_n553), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n740), .A2(new_n744), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n751), .B2(new_n694), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n747), .A2(new_n744), .A3(new_n739), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n612), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n700), .A2(new_n756), .A3(new_n681), .A4(new_n702), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n735), .B1(new_n758), .B2(G330), .ZN(new_n759));
  AOI211_X1 g0559(.A(KEYINPUT87), .B(new_n698), .C1(new_n755), .C2(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n734), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT89), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n734), .A2(KEYINPUT89), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n719), .B1(new_n766), .B2(G1), .ZN(G364));
  INV_X1    g0567(.A(new_n699), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n248), .B1(new_n684), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n714), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n697), .A2(new_n698), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OR3_X1    g0574(.A1(KEYINPUT91), .A2(G13), .A3(G33), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT91), .B1(G13), .B2(G33), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT97), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n697), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n259), .B1(G20), .B2(new_n338), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n540), .A2(new_n713), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n242), .A2(new_n492), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(new_n492), .C2(new_n209), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n255), .A2(new_n213), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n206), .A2(new_n788), .B1(G116), .B2(new_n213), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT90), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n783), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n371), .A2(new_n455), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT93), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n286), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n381), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT95), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT95), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G107), .ZN(new_n800));
  NAND2_X1  g0600(.A1(G20), .A2(G179), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT92), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n381), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n303), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n417), .A2(new_n805), .B1(new_n808), .B2(new_n414), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G20), .A3(new_n381), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(G190), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G20), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n803), .A2(new_n303), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n814), .B1(new_n220), .B2(new_n817), .C1(new_n819), .C2(new_n333), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n794), .A2(G190), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n255), .B1(new_n821), .B2(new_n218), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n809), .B(new_n820), .C1(new_n822), .C2(KEYINPUT94), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n800), .B(new_n823), .C1(KEYINPUT94), .C2(new_n822), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n806), .A2(G200), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(G77), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  INV_X1    g0627(.A(new_n821), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n255), .B1(new_n828), .B2(G303), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n798), .A2(new_n827), .B1(new_n829), .B2(KEYINPUT96), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT96), .ZN(new_n831));
  INV_X1    g0631(.A(new_n811), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n818), .A2(G326), .B1(G329), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  INV_X1    g0634(.A(new_n825), .ZN(new_n835));
  INV_X1    g0635(.A(G322), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n834), .A2(new_n835), .B1(new_n805), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT33), .B(G317), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n807), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n831), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n830), .B(new_n840), .C1(G294), .C2(new_n816), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n782), .B1(new_n826), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n781), .A2(new_n791), .A3(new_n842), .A4(new_n771), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n774), .A2(new_n843), .ZN(G396));
  INV_X1    g0644(.A(new_n761), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n360), .A2(new_n694), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n369), .A2(new_n846), .A3(new_n374), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n369), .A2(new_n846), .A3(new_n374), .A4(KEYINPUT99), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR3_X1    g0651(.A1(new_n369), .A2(KEYINPUT100), .A3(new_n702), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT100), .B1(new_n369), .B2(new_n702), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n722), .A2(new_n723), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n702), .B(new_n855), .C1(new_n662), .C2(new_n670), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n845), .A2(KEYINPUT101), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n858), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n761), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n772), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n761), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n859), .A2(new_n862), .A3(new_n866), .A4(new_n772), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n799), .A2(G87), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n825), .A2(G116), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n828), .A2(G107), .ZN(new_n871));
  INV_X1    g0671(.A(G303), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n827), .A2(new_n808), .B1(new_n819), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G294), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n805), .A2(new_n874), .B1(new_n220), .B2(new_n817), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n314), .B1(new_n811), .B2(new_n834), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n799), .A2(G68), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n540), .B1(new_n817), .B2(new_n417), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n828), .B2(G50), .ZN(new_n881));
  INV_X1    g0681(.A(G132), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n879), .B(new_n881), .C1(new_n882), .C2(new_n811), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT98), .Z(new_n884));
  AOI22_X1  g0684(.A1(G143), .A2(new_n804), .B1(new_n807), .B2(G150), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n885), .B1(new_n886), .B2(new_n819), .C1(new_n812), .C2(new_n835), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT34), .Z(new_n888));
  OAI21_X1  g0688(.A(new_n878), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n772), .B1(new_n889), .B2(new_n782), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n777), .A2(new_n782), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n226), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n778), .C2(new_n855), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n868), .A2(new_n893), .ZN(G384));
  NAND2_X1  g0694(.A1(new_n299), .A2(new_n694), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n300), .A2(new_n309), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n300), .B2(new_n309), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n855), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n752), .B1(new_n651), .B2(new_n702), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n692), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n438), .A2(KEYINPUT16), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n452), .B1(new_n903), .B2(new_n439), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n458), .A2(new_n462), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n902), .B(new_n905), .C1(new_n906), .C2(new_n677), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n461), .A2(new_n902), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n908), .B(new_n431), .C1(new_n909), .C2(new_n453), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n457), .A2(new_n692), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n905), .A2(new_n911), .B1(new_n453), .B2(new_n405), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n908), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n907), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n901), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n459), .B(new_n902), .C1(new_n906), .C2(new_n677), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n431), .B1(new_n909), .B2(new_n453), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n910), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n901), .B(KEYINPUT40), .C1(new_n914), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n751), .A2(new_n694), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT31), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n757), .A2(new_n928), .A3(new_n900), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n465), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n925), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(G330), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n465), .B1(new_n724), .B2(new_n733), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n679), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n914), .B2(new_n923), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n692), .B(new_n904), .C1(new_n450), .C2(new_n463), .ZN(new_n938));
  INV_X1    g0738(.A(new_n913), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(KEYINPUT39), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n300), .A2(new_n694), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n906), .A2(new_n692), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n896), .A2(new_n897), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n369), .A2(new_n694), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n858), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n914), .B2(new_n915), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n934), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n932), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n248), .B2(new_n684), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT35), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n286), .B(new_n259), .C1(new_n535), .C2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(G116), .C1(new_n955), .C2(new_n535), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n717), .A2(new_n226), .A3(new_n418), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n201), .A2(new_n414), .ZN(new_n960));
  OAI211_X1 g0760(.A(G1), .B(new_n683), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(G367));
  OAI211_X1 g0762(.A(new_n564), .B(new_n574), .C1(new_n571), .C2(new_n702), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n667), .A2(new_n694), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n707), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT106), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n709), .A2(new_n963), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n564), .B1(new_n963), .B2(new_n513), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n702), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT103), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n657), .A2(new_n659), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n730), .B1(new_n975), .B2(new_n702), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n975), .A2(new_n611), .A3(new_n702), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n974), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT105), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n973), .A2(new_n985), .A3(new_n981), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n973), .B2(new_n981), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n966), .A2(new_n967), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n968), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n967), .A3(new_n966), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n714), .B(new_n994), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT109), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n709), .B1(new_n513), .B2(new_n694), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(new_n965), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n999), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n965), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n997), .B(new_n707), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n707), .A2(new_n997), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n999), .B(new_n1000), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1003), .B(KEYINPUT44), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n699), .A2(KEYINPUT109), .A3(new_n706), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n699), .B(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n766), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n996), .B1(new_n1014), .B2(new_n766), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n992), .B(new_n993), .C1(new_n1015), .C2(new_n770), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n783), .B1(new_n213), .B2(new_n609), .C1(new_n785), .C2(new_n238), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n980), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n772), .B1(new_n1018), .B2(new_n780), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n799), .A2(G97), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n832), .A2(G317), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n426), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT110), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n828), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT46), .B1(new_n828), .B2(G116), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n835), .A2(new_n827), .B1(new_n469), .B2(new_n817), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n874), .A2(new_n808), .B1(new_n819), .B2(new_n834), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1023), .B(new_n1028), .C1(new_n872), .C2(new_n805), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n799), .A2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n818), .A2(G143), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n314), .B1(new_n832), .B2(G137), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n816), .A2(G68), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n805), .C2(new_n330), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n201), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n812), .A2(new_n808), .B1(new_n835), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n828), .C2(G58), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1030), .A2(new_n1031), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1029), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT47), .Z(new_n1040));
  INV_X1    g0840(.A(new_n782), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1017), .B(new_n1019), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1016), .A2(new_n1042), .ZN(G387));
  OR2_X1    g0843(.A1(new_n766), .A2(new_n1013), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n766), .A2(new_n1013), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n714), .A3(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n712), .B(new_n492), .C1(new_n414), .C2(new_n226), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n327), .A2(new_n333), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1047), .A2(KEYINPUT112), .B1(KEYINPUT50), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT112), .B2(new_n1047), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1048), .A2(KEYINPUT50), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n784), .B1(new_n492), .B2(new_n235), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(G107), .B2(new_n213), .C1(new_n712), .C2(new_n788), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n783), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n706), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n772), .B1(new_n1055), .B2(new_n780), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G311), .A2(new_n807), .B1(new_n804), .B2(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n872), .B2(new_n835), .C1(new_n836), .C2(new_n819), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT48), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n827), .B2(new_n817), .C1(new_n874), .C2(new_n821), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT114), .Z(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n832), .A2(G326), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n540), .B1(new_n799), .B2(G116), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n426), .B1(G150), .B2(new_n832), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n582), .A2(new_n816), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n835), .C2(new_n414), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n333), .A2(new_n805), .B1(new_n819), .B2(new_n812), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n327), .C2(new_n807), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n828), .A2(G77), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1020), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT113), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1054), .B(new_n1056), .C1(new_n1075), .C2(new_n1041), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1013), .A2(new_n770), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT111), .Z(new_n1078));
  NAND3_X1  g0878(.A1(new_n1046), .A2(new_n1076), .A3(new_n1078), .ZN(G393));
  AOI22_X1  g0879(.A1(G150), .A2(new_n818), .B1(new_n804), .B2(G159), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  INV_X1    g0881(.A(new_n327), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1081), .B1(new_n1035), .B2(new_n808), .C1(new_n1082), .C2(new_n835), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n426), .B1(G143), .B2(new_n832), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n869), .B(new_n1084), .C1(new_n414), .C2(new_n821), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT115), .Z(new_n1086));
  AOI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(G77), .C2(new_n816), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G311), .A2(new_n804), .B1(new_n818), .B2(G317), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n828), .B2(G283), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n255), .B1(new_n816), .B2(G116), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n835), .B2(new_n874), .C1(new_n872), .C2(new_n808), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1088), .B2(KEYINPUT52), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n800), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G322), .B2(new_n832), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n782), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n771), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n779), .B2(new_n965), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n783), .B1(new_n220), .B2(new_n213), .C1(new_n785), .C2(new_n245), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n770), .B2(new_n1011), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1011), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1045), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n714), .A3(new_n1014), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(G390));
  NAND3_X1  g0904(.A1(new_n929), .A2(G330), .A3(new_n855), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n946), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n858), .A2(new_n948), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n946), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n943), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n936), .A2(new_n942), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n914), .B2(new_n923), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n732), .A2(new_n702), .A3(new_n855), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n946), .B1(new_n1114), .B2(new_n948), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n914), .A2(new_n915), .A3(new_n935), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n453), .B(new_n692), .C1(new_n450), .C2(new_n463), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n922), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n937), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT39), .B1(new_n1121), .B2(new_n941), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1118), .A2(new_n1122), .B1(new_n943), .B2(new_n949), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n943), .B1(new_n1121), .B2(new_n941), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1114), .A2(new_n948), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n946), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n855), .B(new_n1109), .C1(new_n759), .C2(new_n760), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1123), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1117), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n769), .ZN(new_n1131));
  INV_X1    g0931(.A(G125), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n255), .B1(new_n1132), .B2(new_n811), .C1(new_n798), .C2(new_n1035), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT116), .Z(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n818), .B1(new_n804), .B2(G132), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT117), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AOI22_X1  g0937(.A1(G137), .A2(new_n807), .B1(new_n825), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n821), .A2(new_n330), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT53), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1136), .B(new_n1141), .C1(new_n1140), .C2(new_n1139), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1134), .B(new_n1142), .C1(new_n812), .C2(new_n817), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n469), .A2(new_n808), .B1(new_n805), .B2(new_n624), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n255), .B1(new_n832), .B2(G294), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n226), .B2(new_n817), .C1(new_n819), .C2(new_n827), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G97), .C2(new_n825), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n879), .B(new_n1147), .C1(new_n218), .C2(new_n821), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n771), .B1(new_n1149), .B2(new_n1041), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n778), .B1(new_n936), .B2(new_n942), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n1082), .C2(new_n891), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1131), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1105), .A2(new_n946), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1127), .A2(new_n1125), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n855), .B1(new_n759), .B2(new_n760), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1106), .B1(new_n1156), .B2(new_n946), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1108), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n930), .A2(G330), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n933), .A2(new_n679), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n714), .B1(new_n1130), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1117), .A2(new_n1129), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1153), .B1(new_n1163), .B2(new_n1166), .ZN(G378));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n951), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n895), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n310), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n300), .A2(new_n309), .A3(new_n895), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1171), .A2(new_n1172), .B1(new_n851), .B2(new_n854), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n929), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n940), .B2(new_n941), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n924), .B(G330), .C1(new_n1175), .C2(KEYINPUT40), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n902), .A2(new_n337), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT56), .Z(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT55), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n674), .B2(new_n340), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n672), .A2(new_n673), .A3(KEYINPUT55), .A4(new_n341), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n673), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n387), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n340), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT55), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n674), .A2(new_n1180), .A3(new_n340), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1178), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1176), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1192), .A2(new_n918), .A3(G330), .A4(new_n924), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1169), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1169), .B1(new_n1193), .B2(new_n1191), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n933), .A2(new_n679), .A3(new_n1160), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1165), .B2(new_n1159), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1168), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1161), .B1(new_n1130), .B2(new_n1162), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n951), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1194), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n1204), .A3(KEYINPUT57), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1205), .A3(new_n714), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n772), .B1(new_n1035), .B2(new_n891), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1192), .A2(new_n778), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n799), .A2(G58), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n807), .A2(G97), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G41), .B1(new_n832), .B2(G283), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n426), .A3(new_n1033), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n469), .A2(new_n805), .B1(new_n819), .B2(new_n624), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n582), .C2(new_n825), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1210), .A2(new_n1072), .A3(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G41), .B1(new_n540), .B2(G33), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n807), .B1(new_n825), .B2(G137), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT118), .Z(new_n1220));
  NAND2_X1  g1020(.A1(new_n804), .A2(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n819), .A2(new_n1132), .B1(new_n330), .B2(new_n817), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n828), .B2(new_n1137), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT119), .Z(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G33), .B1(new_n832), .B2(G124), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n263), .B(new_n1228), .C1(new_n798), .C2(new_n812), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT120), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1227), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1217), .B1(G50), .B2(new_n1218), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1208), .B(new_n1209), .C1(new_n782), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1204), .B2(new_n770), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1206), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n825), .A2(G150), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n828), .A2(G159), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n807), .A2(new_n1137), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n805), .B2(new_n886), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n540), .B1(new_n333), .B2(new_n817), .C1(new_n819), .C2(new_n882), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G128), .C2(new_n832), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1210), .A2(new_n1238), .A3(new_n1239), .A4(new_n1243), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n469), .A2(new_n835), .B1(new_n805), .B2(new_n827), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1068), .B1(new_n819), .B2(new_n874), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n314), .B1(new_n811), .B2(new_n872), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1030), .B(new_n1248), .C1(new_n220), .C2(new_n821), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n808), .A2(new_n624), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1244), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n772), .B1(new_n1251), .B2(new_n782), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1109), .B2(new_n778), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n414), .B2(new_n891), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1159), .B2(new_n770), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n995), .B(KEYINPUT122), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1162), .A2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1255), .B1(new_n1257), .B2(new_n1258), .ZN(G381));
  NAND4_X1  g1059(.A1(new_n1016), .A2(new_n1042), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G381), .A2(G384), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1260), .A2(G396), .A3(G393), .A4(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G375), .A2(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(G407));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1262), .B2(new_n693), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G213), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(KEYINPUT60), .A3(new_n1198), .A4(new_n1155), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1273), .A3(new_n714), .A4(new_n1162), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1255), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n893), .A3(new_n868), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G384), .A2(new_n1255), .A3(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1201), .A2(new_n1204), .A3(new_n1256), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1201), .A2(new_n1204), .A3(KEYINPUT123), .A4(new_n1256), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1236), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1206), .A2(G378), .A3(new_n1236), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1269), .B(new_n1278), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1267), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1269), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1278), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1288), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1289), .A2(new_n1290), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1269), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1278), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1276), .A2(new_n1277), .A3(new_n1298), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1292), .B2(new_n1291), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G387), .A2(G390), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1260), .ZN(new_n1307));
  XOR2_X1   g1107(.A(G393), .B(G396), .Z(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(G396), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1306), .A3(new_n1260), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(KEYINPUT63), .B2(new_n1287), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1294), .B1(new_n1303), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1315), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(new_n1314), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1312), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1297), .B2(new_n1304), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1315), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(G405));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1321), .B1(new_n1326), .B2(new_n1293), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1312), .A2(KEYINPUT127), .A3(new_n1278), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1284), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1330), .B(new_n1286), .C1(KEYINPUT127), .C2(new_n1278), .ZN(new_n1331));
  XOR2_X1   g1131(.A(new_n1329), .B(new_n1331), .Z(G402));
endmodule


