//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n213), .A2(new_n214), .B1(new_n205), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n212), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  AND2_X1   g0031(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n233), .A2(new_n210), .A3(new_n234), .ZN(new_n235));
  NOR4_X1   g0035(.A1(new_n228), .A2(new_n231), .A3(new_n232), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  OAI21_X1  g0051(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  AND4_X1   g0061(.A1(new_n255), .A2(new_n259), .A3(new_n261), .A4(G1698), .ZN(new_n262));
  OAI21_X1  g0062(.A(G223), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n261), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n266), .C1(new_n223), .C2(new_n256), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n260), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n254), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n252), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G226), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G190), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n234), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n209), .A2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G50), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n203), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(KEYINPUT8), .A2(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT8), .A2(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n210), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n285), .B1(new_n286), .B2(new_n288), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n284), .B1(new_n295), .B2(new_n280), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n278), .A2(new_n202), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n271), .A2(new_n274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(KEYINPUT9), .A3(new_n297), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n276), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n259), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n256), .A2(KEYINPUT69), .A3(G232), .A4(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n256), .A2(G226), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n254), .B1(new_n315), .B2(new_n270), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n273), .A2(G238), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n316), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g0122(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G179), .A3(new_n320), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(G169), .C1(new_n321), .C2(new_n322), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n288), .A2(new_n202), .B1(new_n294), .B2(new_n223), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n210), .A2(G68), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n280), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT11), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT68), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n277), .B(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n280), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n282), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT12), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G68), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n278), .A2(KEYINPUT12), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n277), .B(KEYINPUT68), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(KEYINPUT12), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n334), .A2(new_n340), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n326), .A2(G190), .A3(new_n320), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n326), .A2(KEYINPUT71), .A3(G190), .A4(new_n320), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  INV_X1    g0152(.A(new_n322), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n320), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n272), .A2(new_n224), .ZN(new_n357));
  OAI21_X1  g0157(.A(G238), .B1(new_n257), .B2(new_n262), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n265), .A2(G232), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n264), .A2(G107), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI211_X1 g0161(.A(new_n254), .B(new_n357), .C1(new_n361), .C2(new_n270), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n270), .ZN(new_n365));
  INV_X1    g0165(.A(new_n254), .ZN(new_n366));
  INV_X1    g0166(.A(new_n357), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n289), .A2(new_n290), .A3(new_n287), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n210), .B2(new_n223), .C1(new_n372), .C2(new_n294), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n280), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n342), .A2(new_n223), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n223), .C2(new_n338), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  AND4_X1   g0177(.A1(new_n307), .A2(new_n346), .A3(new_n356), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT79), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT78), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n260), .A2(new_n213), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT72), .B1(new_n258), .B2(G33), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(G226), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(G1698), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n381), .B(new_n382), .C1(new_n387), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n384), .A2(new_n386), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(new_n390), .A3(new_n259), .ZN(new_n393));
  INV_X1    g0193(.A(new_n382), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT75), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n270), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  INV_X1    g0197(.A(G232), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT76), .B1(new_n272), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n269), .A2(new_n400), .A3(G232), .A4(new_n252), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n254), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n396), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n380), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n393), .A2(new_n394), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n381), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n393), .A2(KEYINPUT75), .A3(new_n394), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n269), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n399), .A2(new_n401), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n366), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n352), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n392), .A2(new_n259), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n210), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT7), .B1(new_n387), .B2(G20), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G68), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G58), .A2(G68), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(G58), .C2(G68), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(G20), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n287), .A2(G159), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT74), .B1(new_n258), .B2(G33), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT74), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n433), .A3(new_n259), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n417), .B1(new_n256), .B2(G20), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n343), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n426), .A2(new_n438), .A3(new_n280), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n293), .B1(new_n209), .B2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n281), .B1(new_n278), .B2(new_n293), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n379), .B1(new_n415), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT79), .B(new_n442), .C1(new_n405), .C2(new_n414), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT17), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n403), .A2(new_n404), .A3(new_n380), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT78), .B1(new_n412), .B2(new_n413), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n442), .B1(new_n405), .B2(new_n414), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT80), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  OAI21_X1  g0257(.A(G169), .B1(new_n409), .B2(new_n411), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n396), .A2(G179), .A3(new_n402), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(new_n442), .A3(KEYINPUT18), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT18), .B1(new_n460), .B2(new_n442), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n442), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT18), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n442), .A3(KEYINPUT18), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(KEYINPUT77), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n275), .A2(new_n363), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n298), .C1(G169), .C2(new_n275), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n365), .A2(G190), .A3(new_n366), .A4(new_n367), .ZN(new_n473));
  INV_X1    g0273(.A(new_n376), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(new_n362), .C2(new_n352), .ZN(new_n475));
  AND4_X1   g0275(.A1(new_n456), .A2(new_n470), .A3(new_n472), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n342), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n209), .B2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n336), .A2(new_n337), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(G20), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n280), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(G33), .B2(G283), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G33), .B2(new_n205), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT20), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n478), .B(new_n480), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n312), .A2(G264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n215), .A2(new_n312), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n387), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT86), .B(G303), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n256), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n269), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n209), .A2(G45), .A3(G274), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n209), .A3(G45), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n499), .A2(G270), .A3(new_n269), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n488), .B1(new_n501), .B2(new_n352), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(G190), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT87), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n488), .B(new_n505), .C1(new_n501), .C2(new_n352), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(G179), .A3(new_n487), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n501), .A2(new_n369), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n487), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n488), .A2(new_n501), .A3(KEYINPUT21), .A4(new_n369), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n507), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n215), .A2(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n214), .A2(new_n312), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n387), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G294), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n269), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n499), .A2(G264), .A3(new_n269), .ZN(new_n520));
  NOR4_X1   g0320(.A1(new_n519), .A2(new_n520), .A3(G179), .A4(new_n498), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n519), .A2(new_n498), .A3(new_n520), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n281), .B1(G1), .B2(new_n260), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n209), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n524), .A2(new_n206), .B1(KEYINPUT25), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n213), .A2(G20), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n387), .A2(KEYINPUT22), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G20), .A3(new_n206), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n260), .A2(new_n477), .A3(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n259), .A3(new_n261), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n528), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n528), .A2(new_n532), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n526), .B1(new_n541), .B2(new_n280), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n525), .A2(KEYINPUT25), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n521), .B(new_n523), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n519), .A2(new_n498), .ZN(new_n545));
  INV_X1    g0345(.A(new_n520), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n522), .A2(G190), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n542), .A2(new_n548), .A3(new_n549), .A4(new_n543), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n514), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n542), .A2(new_n543), .ZN(new_n553));
  INV_X1    g0353(.A(new_n521), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(G169), .C2(new_n522), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n550), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n513), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n277), .A2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n207), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  INV_X1    g0363(.A(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(new_n207), .A3(new_n565), .A4(new_n559), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g0368(.A(G20), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n435), .A2(new_n436), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n287), .A2(G77), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n558), .B1(new_n573), .B2(new_n280), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n524), .A2(new_n205), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n387), .A2(G244), .A3(new_n312), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n312), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT83), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(G33), .B2(G283), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n265), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(G244), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n270), .ZN(new_n587));
  INV_X1    g0387(.A(new_n498), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n499), .A2(G257), .A3(new_n269), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n369), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n577), .B(new_n591), .C1(G179), .C2(new_n590), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n587), .A2(G190), .A3(new_n588), .A4(new_n589), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n574), .A3(new_n576), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n498), .B1(new_n586), .B2(new_n270), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n352), .B1(new_n595), .B2(new_n589), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT84), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n596), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n558), .B(new_n575), .C1(new_n573), .C2(new_n280), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n593), .ZN(new_n601));
  INV_X1    g0401(.A(G45), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n269), .B(G250), .C1(G1), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G238), .A2(G1698), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n224), .B2(G1698), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n387), .A2(new_n605), .B1(G33), .B2(G116), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n496), .B(new_n603), .C1(new_n606), .C2(new_n269), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G190), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n213), .A2(new_n205), .A3(new_n206), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n314), .A2(new_n210), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT19), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n294), .B2(new_n205), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n387), .A2(new_n210), .A3(G68), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n337), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n524), .A2(new_n213), .ZN(new_n618));
  INV_X1    g0418(.A(new_n372), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n336), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n607), .A2(G200), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n609), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n617), .A2(new_n620), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n524), .A2(new_n372), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT85), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n617), .A2(new_n626), .A3(new_n629), .A4(new_n620), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n607), .A2(new_n363), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n607), .A2(G169), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n624), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n592), .A2(new_n597), .A3(new_n601), .A4(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n378), .A2(new_n476), .A3(new_n557), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n472), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT90), .B1(new_n305), .B2(new_n306), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT90), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n461), .A2(new_n462), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT79), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n453), .A2(new_n379), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n649), .A2(KEYINPUT17), .B1(new_n452), .B2(new_n454), .ZN(new_n650));
  INV_X1    g0450(.A(new_n377), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n356), .A2(new_n651), .B1(new_n345), .B2(new_n330), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n639), .B1(new_n643), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n476), .A2(new_n378), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n633), .A2(new_n634), .B1(new_n625), .B2(new_n627), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n624), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n550), .B(new_n657), .C1(new_n658), .C2(new_n544), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n597), .A2(new_n601), .A3(new_n592), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n631), .A2(new_n635), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n623), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n663), .B2(new_n592), .ZN(new_n664));
  INV_X1    g0464(.A(new_n656), .ZN(new_n665));
  INV_X1    g0465(.A(new_n590), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n599), .B1(new_n363), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n657), .A3(new_n668), .A4(new_n591), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n661), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n654), .B1(new_n655), .B2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(G13), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G20), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n209), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n678), .A3(G213), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT91), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n676), .A2(new_n678), .A3(new_n681), .A4(G213), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n488), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n658), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n513), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n552), .A2(new_n556), .B1(new_n553), .B2(new_n685), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n555), .A2(new_n686), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n552), .A2(new_n556), .A3(new_n555), .ZN(new_n695));
  INV_X1    g0495(.A(new_n658), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n555), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n697), .A3(new_n686), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0500(.A(new_n229), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n610), .A2(G116), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n702), .A2(new_n704), .A3(new_n209), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  INV_X1    g0508(.A(new_n702), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n708), .C1(new_n233), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n686), .B1(new_n661), .B2(new_n670), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n665), .A2(new_n623), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n592), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n636), .A2(new_n667), .A3(new_n668), .A4(new_n591), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n665), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n686), .C1(new_n661), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n590), .A2(new_n547), .ZN(new_n721));
  AOI21_X1  g0521(.A(G179), .B1(new_n721), .B2(KEYINPUT95), .ZN(new_n722));
  INV_X1    g0522(.A(new_n501), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n590), .A2(new_n724), .A3(new_n547), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n607), .A4(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n494), .A2(new_n500), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n522), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n666), .A2(new_n729), .A3(KEYINPUT30), .A4(new_n632), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n595), .A2(new_n589), .A3(new_n632), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n728), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n686), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(KEYINPUT31), .B2(new_n735), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n557), .A2(new_n637), .A3(new_n686), .ZN(new_n739));
  OAI21_X1  g0539(.A(G330), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n720), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n711), .B1(new_n741), .B2(G1), .ZN(G364));
  AOI21_X1  g0542(.A(new_n209), .B1(new_n674), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n702), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n689), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n229), .A2(new_n256), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(G87), .B2(new_n207), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n229), .A2(G116), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n701), .A2(new_n387), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n233), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n602), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n247), .A2(G45), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n749), .B(new_n750), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n673), .A2(new_n260), .A3(KEYINPUT96), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G13), .B2(G33), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n234), .B1(G20), .B2(new_n369), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n745), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT97), .Z(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(new_n363), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G58), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n771), .A2(new_n772), .B1(new_n774), .B2(new_n223), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n769), .A2(new_n352), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n397), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n210), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n202), .B1(new_n205), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n768), .A2(new_n397), .A3(G200), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT99), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT99), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n775), .B(new_n780), .C1(G68), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n210), .A2(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n786), .A2(new_n397), .A3(G200), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n256), .B1(new_n787), .B2(new_n213), .C1(new_n206), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n773), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n785), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n264), .B1(new_n787), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n771), .A2(new_n798), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n797), .B(new_n800), .C1(G329), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n779), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G294), .A2(new_n803), .B1(new_n776), .B2(G326), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  INV_X1    g0605(.A(new_n784), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  OAI211_X1 g0607(.A(new_n802), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n774), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n795), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n763), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n762), .B(KEYINPUT101), .Z(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n767), .B(new_n812), .C1(new_n689), .C2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n747), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n376), .A2(new_n685), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT103), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT103), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n376), .A2(new_n685), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n474), .B1(new_n362), .B2(new_n363), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n822), .A2(new_n475), .B1(new_n823), .B2(new_n370), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n370), .A3(new_n686), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT104), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT104), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n819), .A2(new_n821), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n368), .A2(G200), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n376), .B1(new_n362), .B2(G190), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n828), .B(new_n825), .C1(new_n832), .C2(new_n651), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n712), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(new_n740), .ZN(new_n837));
  INV_X1    g0637(.A(new_n745), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n774), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n770), .A2(G143), .B1(new_n840), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n842), .B2(new_n777), .C1(new_n806), .C2(new_n286), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT34), .ZN(new_n844));
  INV_X1    g0644(.A(new_n788), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G68), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n202), .B2(new_n787), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n416), .B(new_n847), .C1(G132), .C2(new_n801), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n844), .B(new_n848), .C1(new_n772), .C2(new_n779), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n774), .A2(new_n477), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n264), .B1(new_n788), .B2(new_n213), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n777), .A2(new_n796), .B1(new_n787), .B2(new_n206), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(G311), .C2(new_n801), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G97), .A2(new_n803), .B1(new_n770), .B2(G294), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT102), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(new_n799), .C2(new_n806), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n849), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n760), .A2(new_n763), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n857), .A2(new_n763), .B1(new_n223), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n859), .B(new_n745), .C1(new_n835), .C2(new_n761), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n839), .A2(new_n860), .ZN(G384));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n443), .A2(new_n683), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n456), .B2(new_n645), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n458), .A2(new_n459), .A3(new_n683), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n442), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(new_n444), .C2(new_n445), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n453), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n862), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n426), .A2(new_n280), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n420), .B2(new_n425), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n441), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n647), .B2(new_n648), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n869), .B1(new_n880), .B2(new_n866), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n469), .B1(new_n446), .B2(new_n455), .ZN(new_n882));
  INV_X1    g0682(.A(new_n683), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n881), .B(KEYINPUT38), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n557), .A2(new_n637), .A3(new_n686), .ZN(new_n887));
  INV_X1    g0687(.A(new_n736), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n735), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n345), .B(new_n354), .C1(new_n349), .C2(new_n350), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n345), .B(new_n685), .C1(new_n891), .C2(new_n330), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n345), .A2(new_n685), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n346), .A2(new_n356), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n834), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT31), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n735), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n884), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n650), .B2(new_n469), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n902), .B2(new_n881), .ZN(new_n903));
  INV_X1    g0703(.A(new_n885), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT106), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n884), .B1(new_n456), .B2(new_n470), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT37), .B1(new_n647), .B2(new_n648), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n878), .B1(new_n444), .B2(new_n445), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n868), .A2(new_n909), .B1(new_n910), .B2(KEYINPUT37), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n862), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n898), .B1(new_n912), .B2(new_n885), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT106), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT40), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n900), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n887), .A2(new_n889), .B1(new_n896), .B2(new_n735), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n655), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n916), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(G330), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n863), .B1(new_n650), .B2(new_n644), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n872), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n922), .B1(new_n924), .B2(new_n904), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n346), .A2(new_n685), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n892), .A2(new_n894), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n825), .B1(new_n712), .B2(new_n834), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n903), .C2(new_n904), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n644), .A2(new_n683), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n714), .A2(new_n476), .A3(new_n378), .A4(new_n719), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n654), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n933), .B(new_n935), .Z(new_n936));
  XNOR2_X1  g0736(.A(new_n921), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n209), .B2(new_n674), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n567), .A2(new_n568), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT35), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n210), .B(new_n234), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(G116), .C1(new_n940), .C2(new_n939), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT105), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT36), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n422), .A2(new_n423), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n753), .A2(G77), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n945), .A2(new_n946), .B1(G50), .B2(new_n343), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n673), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n938), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT107), .Z(G367));
  NOR2_X1   g0750(.A1(new_n599), .A2(new_n686), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n660), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n592), .B2(new_n686), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n552), .A2(new_n556), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n696), .A2(new_n685), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n592), .B1(new_n952), .B2(new_n555), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n686), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n621), .A2(new_n686), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n656), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n715), .B2(new_n961), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n958), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  INV_X1    g0766(.A(KEYINPUT108), .ZN(new_n967));
  INV_X1    g0767(.A(new_n694), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n953), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(KEYINPUT108), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n702), .B(KEYINPUT41), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n953), .A2(new_n698), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n695), .A2(new_n660), .A3(new_n697), .A4(new_n686), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n968), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n692), .A2(new_n693), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n690), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n694), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n955), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n741), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n975), .B1(new_n988), .B2(new_n741), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n972), .B(new_n973), .C1(new_n989), .C2(new_n744), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n779), .A2(new_n343), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G143), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n223), .B2(new_n788), .C1(new_n993), .C2(new_n777), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n772), .A2(new_n787), .B1(new_n774), .B2(new_n202), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n256), .B1(new_n771), .B2(new_n286), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n842), .B2(new_n791), .C1(new_n792), .C2(new_n806), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n771), .A2(new_n492), .B1(new_n774), .B2(new_n799), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G311), .B2(new_n776), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n784), .A2(G294), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n788), .A2(new_n205), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n416), .B1(new_n1004), .B2(new_n791), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G107), .B2(new_n803), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n787), .A2(new_n477), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n998), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT109), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n838), .B1(new_n1012), .B2(new_n763), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n764), .B1(new_n229), .B2(new_n372), .C1(new_n752), .C2(new_n243), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n814), .C2(new_n963), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n985), .A2(new_n744), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n751), .B1(new_n240), .B2(new_n602), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n703), .B2(new_n748), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n343), .A2(new_n223), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n291), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n202), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n704), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n602), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1019), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n701), .A2(new_n206), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n765), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n770), .B1(new_n776), .B2(G322), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n492), .B2(new_n774), .C1(new_n806), .C2(new_n809), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  INV_X1    g0831(.A(G294), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n799), .B2(new_n779), .C1(new_n1032), .C2(new_n787), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n801), .A2(G326), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n387), .B1(new_n845), .B2(G116), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n293), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1041), .A2(new_n784), .B1(G68), .B2(new_n840), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT112), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n803), .A2(new_n619), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n787), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(G77), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n286), .B2(new_n791), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT111), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n771), .A2(new_n202), .B1(new_n777), .B2(new_n792), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1049), .A2(new_n416), .A3(new_n1002), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1040), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1028), .B1(new_n1052), .B2(new_n763), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n982), .A2(new_n813), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n745), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n702), .B1(new_n985), .B2(new_n741), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1017), .B(new_n1055), .C1(new_n987), .C2(new_n1056), .ZN(G393));
  INV_X1    g0857(.A(new_n981), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n986), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n988), .A2(new_n1059), .A3(new_n702), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n981), .A2(new_n744), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n387), .B1(new_n993), .B2(new_n791), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n803), .A2(G77), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n343), .B2(new_n787), .C1(new_n213), .C2(new_n788), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(new_n1021), .C2(new_n840), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n776), .B1(new_n770), .B2(G159), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n202), .C2(new_n806), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT114), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n779), .A2(new_n477), .B1(new_n774), .B2(new_n1032), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n264), .B1(new_n791), .B2(new_n798), .C1(new_n206), .C2(new_n788), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G283), .C2(new_n1045), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n492), .B2(new_n806), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n770), .B1(new_n776), .B2(G317), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n838), .B1(new_n1076), .B2(new_n763), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n764), .B1(new_n205), .B2(new_n229), .C1(new_n752), .C2(new_n250), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n762), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n1078), .C1(new_n953), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1060), .A2(new_n1061), .A3(new_n1080), .ZN(G390));
  AND3_X1   g0881(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT39), .B1(new_n874), .B2(new_n885), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n760), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n801), .A2(G294), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1063), .A2(new_n264), .A3(new_n846), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G116), .A2(new_n770), .B1(new_n776), .B2(G283), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n213), .B2(new_n787), .C1(new_n205), .C2(new_n774), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G107), .C2(new_n784), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n845), .A2(G50), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n264), .B1(new_n770), .B2(G132), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n801), .A2(G125), .ZN(new_n1092));
  OR3_X1    g0892(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n286), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT53), .B1(new_n787), .B2(new_n286), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G159), .A2(new_n803), .B1(new_n776), .B2(G128), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n774), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1095), .B(new_n1099), .C1(G137), .C2(new_n784), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1089), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT117), .Z(new_n1102));
  AOI21_X1  g0902(.A(new_n838), .B1(new_n1102), .B2(new_n763), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n858), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1084), .B(new_n1103), .C1(new_n1041), .C2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n827), .A2(new_n833), .A3(G330), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n917), .A2(new_n929), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n926), .B1(new_n930), .B2(new_n929), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n925), .B2(new_n927), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n926), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n686), .B1(new_n661), .B2(new_n718), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n825), .B1(new_n1112), .B2(new_n834), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n929), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n892), .A2(KEYINPUT115), .A3(new_n894), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n886), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1108), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1109), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n929), .B(new_n1107), .C1(new_n738), .C2(new_n739), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1119), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1105), .B1(new_n1128), .B2(new_n743), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n917), .A2(new_n476), .A3(new_n378), .A4(G330), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n654), .A2(new_n934), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n661), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n716), .A2(new_n717), .A3(new_n665), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n685), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n826), .B1(new_n1134), .B2(new_n835), .ZN(new_n1135));
  AOI221_X4 g0935(.A(new_n1106), .B1(new_n896), .B2(new_n735), .C1(new_n887), .C2(new_n889), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1124), .B(new_n1135), .C1(new_n1136), .C2(new_n1117), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n930), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1107), .B1(new_n738), .B2(new_n739), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n929), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n1108), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1131), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1110), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1108), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1123), .B2(new_n1119), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT116), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT116), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1127), .A2(new_n1151), .A3(new_n1145), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1150), .A2(new_n1152), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1129), .B1(new_n1153), .B2(new_n702), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G378));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n298), .A2(new_n883), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT56), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n641), .A2(new_n472), .A3(new_n642), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT55), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(KEYINPUT55), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1159), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT55), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n643), .A2(new_n1166), .A3(new_n472), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1161), .A3(new_n1158), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n933), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(new_n928), .A3(new_n931), .A4(new_n932), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n900), .C1(new_n907), .C2(new_n915), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT118), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1170), .A2(new_n1174), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1131), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n709), .B1(new_n1182), .B2(KEYINPUT57), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1131), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT119), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1151), .B1(new_n1127), .B2(new_n1145), .ZN(new_n1189));
  AOI211_X1 g0989(.A(KEYINPUT116), .B(new_n1144), .C1(new_n1121), .C2(new_n1126), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1131), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AND4_X1   g0991(.A1(new_n1170), .A2(new_n1174), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1170), .A2(new_n1172), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1184), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1183), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1194), .A2(new_n744), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n801), .A2(G283), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n992), .A2(new_n268), .A3(new_n1046), .A4(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n771), .A2(new_n206), .B1(new_n777), .B2(new_n477), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n788), .A2(new_n772), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n774), .A2(new_n372), .ZN(new_n1204));
  OR4_X1    g1004(.A1(new_n387), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1201), .B(new_n1205), .C1(G97), .C2(new_n784), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  NAND2_X1  g1007(.A1(new_n784), .A2(G132), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n770), .A2(G128), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n776), .A2(G125), .B1(new_n840), .B2(G137), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n803), .A2(G150), .B1(new_n1045), .B2(new_n1097), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT59), .Z(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n845), .B2(G159), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G33), .B1(new_n801), .B2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G41), .B1(new_n387), .B2(G33), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1207), .B(new_n1216), .C1(G50), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n838), .B1(new_n1218), .B2(new_n763), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(G50), .B2(new_n1104), .C1(new_n1175), .C2(new_n761), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1199), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1156), .B1(new_n1198), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1198), .A2(new_n1156), .A3(new_n1221), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(G375));
  NOR2_X1   g1025(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(new_n743), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1115), .A2(new_n760), .A3(new_n1116), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT121), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n787), .A2(new_n792), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n779), .A2(new_n202), .B1(new_n774), .B2(new_n286), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G137), .C2(new_n770), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n776), .A2(G132), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n784), .A2(new_n1097), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n416), .B(new_n1203), .C1(G128), .C2(new_n801), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n264), .B1(new_n788), .B2(new_n223), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1044), .B1(new_n206), .B2(new_n774), .C1(new_n777), .C2(new_n1032), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G283), .C2(new_n770), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n477), .B2(new_n806), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n787), .A2(new_n205), .B1(new_n791), .B2(new_n796), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT122), .Z(new_n1243));
  OAI21_X1  g1043(.A(new_n1237), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1244), .A2(new_n763), .B1(new_n343), .B2(new_n858), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1229), .A2(new_n1230), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1227), .B1(new_n745), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1226), .A2(new_n1185), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n974), .A3(new_n1144), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(G381));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n990), .A2(new_n1015), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G381), .A2(G384), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT123), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1198), .A2(new_n1156), .A3(new_n1221), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n1222), .A3(G378), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1253), .A2(KEYINPUT123), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1258), .A2(new_n1260), .A3(KEYINPUT124), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1223), .A2(new_n1154), .A3(new_n1224), .A4(new_n1261), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1257), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(G407));
  NAND3_X1  g1066(.A1(new_n1223), .A2(new_n1154), .A3(new_n1224), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G343), .C2(new_n1267), .ZN(G409));
  AOI21_X1  g1068(.A(new_n1154), .B1(new_n1198), .B2(new_n1221), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n702), .B(new_n1144), .C1(new_n1248), .C2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT60), .B1(new_n1226), .B2(new_n1185), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1247), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n839), .A3(new_n860), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1247), .B(G384), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1182), .A2(new_n974), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1221), .A2(new_n1277), .A3(new_n1154), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n684), .A2(G213), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1269), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1221), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1196), .B1(new_n1195), .B2(new_n1184), .ZN(new_n1287));
  AOI211_X1 g1087(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n1191), .C2(new_n1194), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1289), .B2(new_n1183), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1284), .B(new_n1285), .C1(new_n1290), .C2(new_n1154), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1284), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1276), .A2(KEYINPUT125), .A3(new_n1293), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1296), .A2(new_n1297), .B1(new_n1295), .B2(new_n1284), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1269), .B2(new_n1280), .ZN(new_n1299));
  XOR2_X1   g1099(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1300));
  NAND4_X1  g1100(.A1(new_n1283), .A2(new_n1292), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(G393), .B(new_n816), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1251), .B1(new_n990), .B2(new_n1015), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1253), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1302), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1252), .A3(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1311), .B(new_n1308), .C1(new_n1281), .C2(KEYINPUT63), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1299), .B2(new_n1291), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1312), .A2(new_n1314), .A3(KEYINPUT126), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1284), .A2(new_n1295), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1191), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n702), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1287), .A2(new_n1288), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(G378), .B1(new_n1322), .B2(new_n1286), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1319), .B1(new_n1323), .B2(new_n1285), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT63), .B1(new_n1324), .B2(new_n1281), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1304), .A2(new_n1311), .A3(new_n1307), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1291), .B2(new_n1313), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1316), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1310), .B1(new_n1315), .B2(new_n1328), .ZN(G405));
  OAI21_X1  g1129(.A(new_n1284), .B1(new_n1260), .B2(new_n1269), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1267), .A2(new_n1276), .A3(new_n1323), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1330), .A2(new_n1308), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1308), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


