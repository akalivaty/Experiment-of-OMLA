//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  XNOR2_X1  g033(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(KEYINPUT68), .B1(G567), .B2(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT69), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT69), .B1(new_n466), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n473), .A2(G2105), .B1(new_n479), .B2(new_n481), .ZN(G160));
  NAND3_X1  g057(.A1(new_n466), .A2(new_n468), .A3(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n466), .A2(new_n468), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n491), .B2(KEYINPUT71), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n485), .B(new_n492), .C1(KEYINPUT71), .C2(new_n491), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n493), .A2(KEYINPUT73), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  AND2_X1   g072(.A1(KEYINPUT74), .A2(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT74), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2105), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n508), .A2(new_n466), .A3(new_n468), .A4(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n467), .A2(G2104), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT4), .B1(new_n519), .B2(new_n508), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n513), .A2(new_n520), .ZN(G164));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT6), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G50), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI221_X1 g113(.A(KEYINPUT76), .B1(new_n534), .B2(new_n535), .C1(new_n533), .C2(new_n532), .ZN(new_n539));
  NAND2_X1  g114(.A1(G75), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(new_n525), .ZN(new_n541));
  INV_X1    g116(.A(G62), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n538), .A2(new_n539), .B1(G651), .B2(new_n543), .ZN(G166));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT77), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT7), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(new_n530), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G89), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n522), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G51), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n547), .A2(new_n554), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  INV_X1    g132(.A(G52), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n532), .A2(new_n557), .B1(new_n534), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n527), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(G171));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n532), .A2(new_n563), .B1(new_n534), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n527), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n551), .A2(G53), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n541), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(G651), .A2(new_n579), .B1(new_n549), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  NAND2_X1  g157(.A1(new_n538), .A2(new_n539), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n543), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n549), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n551), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n541), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(KEYINPUT78), .A3(G651), .ZN(new_n596));
  AOI22_X1  g171(.A1(G86), .A2(new_n549), .B1(new_n551), .B2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n532), .A2(new_n599), .B1(new_n534), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n527), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n551), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n527), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT79), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n549), .A2(G92), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT10), .Z(new_n612));
  AND2_X1   g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(G299), .B(KEYINPUT80), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n519), .A2(new_n476), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n484), .A2(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT82), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n633), .A2(KEYINPUT82), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n490), .A2(G135), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n630), .A2(new_n631), .A3(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT16), .B(G1341), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n646), .B2(new_n652), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n662), .A2(KEYINPUT17), .A3(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n662), .B2(KEYINPUT17), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n663), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n672), .A2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1991), .ZN(new_n685));
  INV_X1    g260(.A(G1996), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n684), .A2(G1991), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(G1991), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(G1996), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n689), .B1(new_n687), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n670), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n669), .A3(new_n693), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G35), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G162), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT29), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G2090), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G160), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n700), .A2(G33), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G103), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(KEYINPUT25), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(KEYINPUT25), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n717), .B(new_n718), .C1(G139), .C2(new_n490), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n519), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n474), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(new_n700), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n713), .B(new_n714), .C1(G2072), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n726), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n700), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n700), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n724), .A2(G2072), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(G2078), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G299), .ZN(new_n738));
  OAI21_X1  g313(.A(KEYINPUT23), .B1(new_n738), .B2(new_n726), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n726), .A2(G20), .ZN(new_n740));
  MUX2_X1   g315(.A(new_n739), .B(KEYINPUT23), .S(new_n740), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n726), .A2(G4), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n613), .B2(new_n726), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT88), .B(G1348), .Z(new_n744));
  OAI22_X1  g319(.A1(new_n741), .A2(G1956), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n741), .A2(G1956), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n638), .A2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G171), .B2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G1961), .ZN(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT30), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G11), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n726), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n568), .B2(new_n726), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n761), .C1(G1961), .C2(new_n750), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n745), .A2(new_n746), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n725), .A2(new_n737), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n700), .A2(G26), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n484), .A2(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n490), .A2(G140), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n474), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n700), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n765), .B(new_n772), .S(KEYINPUT28), .Z(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2067), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(G2067), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n743), .C2(new_n744), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n700), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n490), .A2(G141), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT26), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n476), .A2(G105), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n484), .A2(G129), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT91), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT91), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n777), .B1(new_n786), .B2(new_n700), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT92), .Z(new_n788));
  XOR2_X1   g363(.A(KEYINPUT27), .B(G1996), .Z(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n776), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n704), .A2(new_n764), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n726), .A2(G24), .ZN(new_n795));
  OAI211_X1 g370(.A(KEYINPUT85), .B(new_n795), .C1(new_n604), .C2(new_n726), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT85), .B2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1986), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n700), .A2(G25), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(G107), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G2105), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n490), .A2(G131), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT84), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n484), .A2(G119), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n799), .B1(new_n808), .B2(new_n700), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G23), .ZN(new_n812));
  XOR2_X1   g387(.A(G288), .B(KEYINPUT86), .Z(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G16), .A2(G22), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G166), .B2(G16), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT87), .B(G1971), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G6), .B(G305), .S(G16), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT32), .B(G1981), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n816), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n798), .B(new_n811), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n794), .A2(new_n831), .ZN(G311));
  OAI21_X1  g407(.A(KEYINPUT95), .B1(new_n794), .B2(new_n831), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n793), .B(new_n834), .C1(new_n829), .C2(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G150));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n532), .A2(new_n837), .B1(new_n534), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n527), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n839), .A2(new_n841), .A3(KEYINPUT96), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT96), .B1(new_n839), .B2(new_n841), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n568), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n842), .B(KEYINPUT96), .C1(new_n567), .C2(new_n565), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n613), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT97), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n845), .B1(new_n859), .B2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n504), .B1(new_n500), .B2(KEYINPUT75), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n511), .B1(new_n863), .B2(new_n503), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n508), .B1(new_n469), .B2(new_n470), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT4), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT100), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n864), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n771), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(new_n786), .ZN(new_n875));
  INV_X1    g450(.A(new_n786), .ZN(new_n876));
  INV_X1    g451(.A(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n872), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n723), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n878), .A3(new_n721), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n862), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n879), .B2(new_n723), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n484), .A2(G130), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n490), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n474), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n886), .B2(KEYINPUT102), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n808), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n808), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n885), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n628), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n628), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n884), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n900), .A2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n882), .B2(new_n883), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n496), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n638), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n884), .B2(new_n904), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n906), .B(KEYINPUT104), .C1(new_n882), .C2(new_n883), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(G395));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  INV_X1    g497(.A(new_n813), .ZN(new_n923));
  NOR2_X1   g498(.A1(G303), .A2(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NOR2_X1   g500(.A1(G166), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n604), .B(G305), .Z(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g504(.A1(G166), .A2(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n813), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n928), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n922), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT108), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n938), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT109), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n623), .B(KEYINPUT105), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(new_n850), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n613), .A2(G299), .ZN(new_n948));
  AOI21_X1  g523(.A(G299), .B1(new_n610), .B2(new_n612), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n850), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n946), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n610), .A2(new_n612), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(new_n738), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(new_n949), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(KEYINPUT41), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n941), .B(new_n963), .C1(KEYINPUT42), .C2(new_n943), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n945), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n945), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G868), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n842), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(G295));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n969), .ZN(G331));
  NAND3_X1  g546(.A1(new_n848), .A2(new_n849), .A3(G301), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G301), .B1(new_n848), .B2(new_n849), .ZN(new_n974));
  OAI21_X1  g549(.A(G286), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n974), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(G168), .A3(new_n972), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n959), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n977), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(new_n960), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n940), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n960), .A2(new_n977), .A3(new_n975), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n939), .B(new_n934), .C1(new_n983), .C2(new_n978), .ZN(new_n984));
  INV_X1    g559(.A(G37), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT110), .B1(new_n959), .B2(new_n955), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  INV_X1    g565(.A(new_n955), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n951), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n959), .A2(KEYINPUT41), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n980), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n978), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n934), .A2(new_n939), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT111), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n981), .B2(new_n940), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n940), .B1(new_n996), .B2(new_n995), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n985), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n988), .B1(new_n1003), .B2(new_n987), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n1003), .B2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(G397));
  XNOR2_X1  g585(.A(new_n771), .B(G2067), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n870), .B2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(G125), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n517), .B2(new_n518), .ZN(new_n1016));
  INV_X1    g591(.A(new_n472), .ZN(new_n1017));
  OAI21_X1  g592(.A(G2105), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n479), .A2(new_n481), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(G40), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1012), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1024));
  INV_X1    g599(.A(new_n808), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(new_n810), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n810), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n786), .B(new_n686), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1024), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1022), .A2(G1986), .A3(G290), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n1021), .B2(new_n686), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1012), .A2(new_n786), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n1021), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1021), .A2(KEYINPUT46), .A3(new_n686), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1038), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1032), .A2(new_n1034), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1024), .A2(new_n1027), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1043));
  INV_X1    g618(.A(G2067), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n771), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1022), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n595), .A2(new_n597), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n596), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(G305), .B2(G1981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G305), .A2(G1981), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT117), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G305), .A2(new_n1056), .A3(G1981), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(KEYINPUT118), .A2(KEYINPUT49), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1053), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1020), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1384), .B1(new_n864), .B2(new_n867), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1060), .B1(new_n1058), .B2(new_n1053), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1065), .A4(new_n1061), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  OR2_X1    g647(.A1(G288), .A2(G1976), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1053), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n813), .A2(G1976), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1065), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1075), .A2(new_n1065), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1082));
  INV_X1    g657(.A(G1384), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT45), .B(new_n1083), .C1(new_n868), .C2(new_n869), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n513), .B2(new_n520), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1020), .B1(new_n1013), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1971), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1020), .B1(KEYINPUT50), .B2(new_n1085), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n1083), .C1(new_n513), .C2(new_n520), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G2090), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G166), .B2(new_n1062), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT115), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G166), .A2(new_n1062), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT114), .B1(new_n1096), .B2(KEYINPUT55), .ZN(new_n1097));
  AND4_X1   g672(.A1(KEYINPUT114), .A2(G303), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g674(.A(G8), .B1(new_n1087), .B2(new_n1092), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1074), .A2(new_n1065), .B1(new_n1082), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1092), .B2(new_n1087), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1064), .A2(KEYINPUT45), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1966), .B1(new_n1086), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1085), .A2(KEYINPUT50), .ZN(new_n1108));
  AND4_X1   g683(.A1(new_n712), .A2(new_n1108), .A3(new_n1063), .A4(new_n1090), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1110), .A2(new_n1062), .A3(G286), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1082), .A2(new_n1100), .A3(new_n1105), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1112), .B2(KEYINPUT120), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1102), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1020), .B2(new_n1085), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1064), .A2(G160), .A3(KEYINPUT121), .A4(G40), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(KEYINPUT122), .A4(new_n1044), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  OAI211_X1 g696(.A(G40), .B(G160), .C1(new_n1064), .C2(new_n1089), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1090), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(new_n1119), .A3(new_n1044), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n957), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n957), .A2(new_n1128), .A3(new_n1124), .A4(new_n1120), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G299), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n576), .A2(new_n580), .A3(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT56), .B(G2072), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1084), .A2(new_n1086), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1956), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1084), .A2(new_n1086), .A3(new_n1137), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1143), .A3(new_n1135), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1128), .A2(new_n1124), .A3(new_n1120), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G1996), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT58), .B(G1341), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n568), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n568), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1144), .A2(KEYINPUT61), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT123), .B1(new_n1160), .B2(new_n1136), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1162), .B(new_n1135), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1159), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1131), .A2(new_n1149), .A3(new_n1158), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1140), .A2(new_n1162), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1160), .A2(KEYINPUT123), .A3(new_n1136), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1128), .A2(new_n1124), .A3(new_n1120), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1167), .A2(new_n1168), .B1(new_n613), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1144), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1173));
  OAI211_X1 g748(.A(KEYINPUT124), .B(new_n1144), .C1(new_n1173), .C2(new_n1129), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1165), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1150), .B2(G2078), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT127), .B(G1961), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1091), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1176), .A2(G2078), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1086), .A2(new_n1106), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G171), .B(KEYINPUT54), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1014), .A2(new_n1063), .A3(new_n1084), .A4(new_n1180), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1177), .A2(new_n1186), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT125), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1189));
  OAI211_X1 g764(.A(G40), .B(G160), .C1(new_n1064), .C2(KEYINPUT45), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1085), .A2(new_n1013), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n729), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1088), .A2(new_n712), .A3(new_n1090), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(G286), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT51), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1197), .A2(new_n1062), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT126), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1194), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1202));
  OAI21_X1  g777(.A(G168), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1203), .A2(new_n1204), .A3(new_n1198), .ZN(new_n1205));
  NOR2_X1   g780(.A1(G168), .A2(new_n1062), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(KEYINPUT51), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1110), .B2(new_n1062), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1200), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1189), .A2(new_n1195), .A3(new_n1206), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1188), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1175), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1209), .A2(new_n1213), .A3(new_n1210), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1182), .A2(G171), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1213), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1212), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AND3_X1   g793(.A1(new_n1082), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1116), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n604), .B(G1986), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1022), .A2(new_n1221), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n1032), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1047), .B1(new_n1220), .B2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g799(.A1(G227), .A2(new_n463), .A3(G401), .ZN(new_n1226));
  AND3_X1   g800(.A1(new_n696), .A2(new_n698), .A3(new_n1226), .ZN(new_n1227));
  AND3_X1   g801(.A1(new_n1227), .A2(new_n917), .A3(new_n1007), .ZN(G308));
  NAND3_X1  g802(.A1(new_n1227), .A2(new_n917), .A3(new_n1007), .ZN(G225));
endmodule


