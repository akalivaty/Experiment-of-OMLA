//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT66), .B(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g0025(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(new_n203), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT65), .Z(new_n234));
  OAI221_X1 g0034(.A(new_n213), .B1(KEYINPUT1), .B2(new_n222), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n248), .B(KEYINPUT68), .Z(new_n249));
  NAND2_X1  g0049(.A1(new_n201), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n226), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(G223), .B1(new_n266), .B2(G77), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n259), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G179), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n204), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n229), .A2(G33), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n283), .B1(new_n284), .B2(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n225), .A2(new_n226), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n289), .A2(new_n291), .B1(new_n201), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n277), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G50), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n270), .A2(new_n280), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(G169), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n282), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n294), .A2(new_n297), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n302), .A2(KEYINPUT9), .B1(new_n281), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n298), .A2(new_n305), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n304), .B2(new_n307), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n268), .A2(G232), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n261), .A2(new_n262), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G238), .A3(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n266), .A2(G107), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n259), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n275), .ZN(new_n321));
  INV_X1    g0121(.A(new_n214), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n274), .A2(new_n278), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n320), .A2(new_n328), .A3(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(new_n291), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT70), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n229), .A3(G33), .ZN(new_n333));
  INV_X1    g0133(.A(new_n287), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G13), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G1), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT71), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n292), .A2(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n330), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n296), .A2(G77), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(G77), .B2(new_n342), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n327), .A2(new_n329), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n320), .A2(G190), .A3(new_n324), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n306), .B1(new_n320), .B2(new_n324), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G232), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G1698), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n312), .B1(G33), .B2(G97), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n357), .A2(new_n259), .B1(new_n321), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT73), .ZN(new_n361));
  INV_X1    g0161(.A(G238), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n275), .A2(KEYINPUT72), .B1(new_n279), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT13), .A4(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(new_n359), .C2(new_n363), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(G169), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT14), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n360), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n360), .B2(new_n364), .ZN(new_n373));
  OAI21_X1  g0173(.A(G179), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT14), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n365), .A2(new_n375), .A3(G169), .A4(new_n368), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT12), .B1(new_n342), .B2(G68), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n203), .A2(G20), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT12), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n338), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n342), .A2(new_n330), .A3(G68), .A4(new_n296), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n201), .A2(KEYINPUT75), .A3(G20), .A4(G33), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n285), .B2(G50), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n379), .B1(new_n288), .B2(new_n215), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n385), .B1(new_n391), .B2(new_n330), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT11), .B(new_n291), .C1(new_n389), .C2(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n384), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n377), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G190), .B1(new_n372), .B2(new_n373), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n365), .A2(G200), .A3(new_n368), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n310), .A2(new_n353), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n261), .A2(new_n229), .A3(new_n262), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n262), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n232), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n285), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n405), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n266), .B2(new_n229), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n264), .A2(new_n265), .A3(new_n407), .A4(G20), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n415), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(new_n424), .A3(new_n291), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n426), .B(new_n427), .ZN(new_n428));
  OR2_X1    g0228(.A1(G223), .A2(G1698), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n276), .A2(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(new_n264), .C2(new_n265), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n318), .ZN(new_n433));
  INV_X1    g0233(.A(G274), .ZN(new_n434));
  INV_X1    g0234(.A(new_n223), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n256), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n323), .A2(G232), .B1(new_n273), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n437), .A3(new_n303), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n259), .B1(new_n428), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n275), .B1(new_n355), .B2(new_n279), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n306), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n287), .B1(new_n277), .B2(G20), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n295), .A2(new_n443), .B1(new_n293), .B2(new_n287), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n425), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT17), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n433), .A2(new_n437), .A3(new_n328), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n326), .B1(new_n439), .B2(new_n440), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n425), .B2(new_n444), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI211_X1 g0252(.A(KEYINPUT18), .B(new_n449), .C1(new_n425), .C2(new_n444), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT79), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  INV_X1    g0255(.A(new_n444), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n422), .A2(new_n423), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n330), .B1(new_n457), .B2(new_n405), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n424), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT18), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n451), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n446), .B1(new_n454), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n404), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n272), .A2(G1), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(G250), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n434), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n274), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G238), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT83), .B1(new_n263), .B2(G244), .ZN(new_n472));
  OAI211_X1 g0272(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(KEYINPUT84), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n318), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n469), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n474), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n312), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n328), .B(new_n468), .C1(new_n477), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G33), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n291), .A2(new_n293), .A3(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT86), .B1(new_n332), .B2(new_n486), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n229), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G87), .B2(new_n208), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n229), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n288), .B2(new_n206), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n330), .B1(new_n496), .B2(KEYINPUT85), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(new_n498), .A3(new_n493), .A4(new_n495), .ZN(new_n499));
  INV_X1    g0299(.A(new_n332), .ZN(new_n500));
  INV_X1    g0300(.A(new_n342), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n497), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n468), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n259), .B1(new_n481), .B2(KEYINPUT84), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n471), .B1(new_n472), .B2(new_n475), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n483), .B(new_n503), .C1(new_n509), .C2(G169), .ZN(new_n510));
  OAI211_X1 g0310(.A(G190), .B(new_n468), .C1(new_n477), .C2(new_n482), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n497), .A2(new_n499), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n500), .A2(new_n501), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n486), .A2(G87), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n511), .B(new_n515), .C1(new_n509), .C2(new_n306), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n277), .B(G45), .C1(new_n271), .C2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT5), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G41), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n274), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT82), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(G41), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n465), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(G257), .A4(new_n274), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT81), .B1(new_n465), .B2(new_n524), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n274), .A2(G274), .A3(new_n523), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n522), .A2(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G283), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n484), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G250), .A2(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT4), .A2(G244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n312), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n318), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n537), .B2(new_n543), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n534), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n550), .A2(new_n206), .A3(G107), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n553), .A2(new_n229), .B1(new_n215), .B2(new_n286), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n207), .B1(new_n408), .B2(new_n409), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n291), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n292), .A2(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n486), .B2(G97), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n534), .B(G190), .C1(new_n546), .C2(new_n547), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n549), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n548), .A2(new_n326), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n534), .B(new_n328), .C1(new_n546), .C2(new_n547), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n558), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT23), .B1(new_n229), .B2(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n207), .A3(G20), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT89), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n229), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n312), .A2(new_n577), .A3(new_n229), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n574), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n291), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n293), .A2(new_n207), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n486), .A2(G107), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n590));
  OAI211_X1 g0390(.A(G250), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n591));
  INV_X1    g0391(.A(G294), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(new_n484), .C2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n525), .A2(new_n274), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n593), .A2(new_n318), .B1(new_n594), .B2(G264), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n518), .A2(new_n528), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n524), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n436), .A3(new_n597), .A4(new_n523), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(G190), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n318), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(G264), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n583), .A2(new_n589), .A3(new_n599), .A4(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n561), .A2(new_n565), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n517), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n607));
  OAI211_X1 g0407(.A(G257), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n261), .A2(G303), .A3(new_n262), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n318), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n525), .A2(G270), .A3(new_n274), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n318), .A3(KEYINPUT87), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n485), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n342), .A2(new_n330), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT88), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(G20), .B1(G33), .B2(G283), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n484), .A2(G97), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n625), .B1(G20), .B2(new_n619), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n291), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n626), .A2(new_n291), .A3(KEYINPUT20), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n501), .A2(new_n619), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n342), .A2(new_n330), .A3(KEYINPUT88), .A4(new_n620), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n623), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n618), .B(new_n635), .C1(new_n303), .C2(new_n617), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n602), .A2(new_n326), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n595), .A2(new_n328), .A3(new_n598), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n574), .A2(new_n579), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT24), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n330), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n637), .B(new_n638), .C1(new_n642), .C2(new_n588), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n634), .A2(new_n617), .A3(G169), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT21), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n634), .A2(new_n617), .A3(KEYINPUT21), .A4(G169), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n617), .A2(new_n328), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n634), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n643), .A2(new_n646), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n464), .A2(new_n606), .A3(new_n636), .A4(new_n651), .ZN(G372));
  NAND2_X1  g0452(.A1(new_n308), .A2(new_n309), .ZN(new_n653));
  INV_X1    g0453(.A(new_n446), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n348), .A2(new_n403), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n400), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n452), .B2(new_n453), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n461), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n653), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n301), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT91), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n404), .A2(new_n463), .ZN(new_n668));
  INV_X1    g0468(.A(new_n510), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n606), .B2(new_n650), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n510), .A3(new_n516), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n510), .A2(new_n671), .A3(new_n516), .A4(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n667), .B1(new_n668), .B2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n646), .A2(new_n649), .A3(new_n647), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n338), .A2(new_n229), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n338), .A2(new_n684), .A3(new_n229), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT92), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT93), .B(G343), .Z(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n681), .A2(new_n636), .B1(new_n634), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n680), .A2(new_n635), .A3(new_n691), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n642), .A2(new_n588), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n604), .B1(new_n698), .B2(new_n691), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(new_n643), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n643), .A2(new_n692), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n681), .A2(new_n692), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(G87), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n206), .A3(new_n207), .A4(new_n619), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT94), .ZN(new_n709));
  INV_X1    g0509(.A(new_n211), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n709), .A2(new_n277), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n233), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  OAI211_X1 g0515(.A(new_n468), .B(new_n595), .C1(new_n477), .C2(new_n482), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n505), .A2(new_n508), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(KEYINPUT96), .A3(new_n468), .A4(new_n595), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n548), .A2(new_n617), .A3(new_n328), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n548), .A2(new_n617), .A3(new_n328), .A4(new_n602), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n509), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n692), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n606), .A2(new_n636), .A3(new_n651), .A4(new_n691), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT31), .ZN(new_n732));
  INV_X1    g0532(.A(G330), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n727), .B1(new_n722), .B2(new_n723), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n691), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n692), .B1(new_n670), .B2(new_n676), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n468), .B1(new_n477), .B2(new_n482), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n744), .A2(new_n326), .B1(new_n502), .B2(new_n489), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n509), .B2(G190), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(G200), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n483), .A2(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n561), .A2(new_n565), .A3(new_n604), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n650), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT98), .ZN(new_n752));
  AND4_X1   g0552(.A1(KEYINPUT26), .A2(new_n671), .A3(new_n510), .A4(new_n516), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n669), .B1(new_n753), .B2(KEYINPUT97), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT97), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n674), .A2(new_n755), .A3(new_n675), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n606), .A2(new_n757), .A3(new_n650), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n752), .A2(new_n754), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n739), .B1(new_n743), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n715), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n710), .A2(new_n266), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n763), .A2(G355), .B1(new_n619), .B2(new_n710), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n710), .A2(new_n312), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n234), .B2(G45), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n254), .A2(new_n272), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT100), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n228), .B1(G20), .B2(new_n326), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n770), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n711), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n337), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n277), .B1(new_n779), .B2(G45), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(KEYINPUT99), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT99), .ZN(new_n782));
  INV_X1    g0582(.A(new_n780), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n711), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n229), .A2(new_n328), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n266), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n787), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(new_n303), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G322), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n229), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n788), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n791), .B(new_n796), .C1(G329), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G326), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n792), .A2(G190), .A3(new_n306), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n804), .A2(new_n805), .B1(G303), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n797), .A2(new_n303), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n328), .A2(new_n306), .A3(G190), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n810), .A2(G283), .B1(new_n812), .B2(G294), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n800), .A2(new_n803), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n806), .A2(new_n707), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n799), .A2(G159), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(KEYINPUT32), .B1(new_n201), .B2(new_n801), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G68), .C2(new_n804), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n812), .B(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G97), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n312), .B1(new_n794), .B2(new_n202), .ZN(new_n821));
  INV_X1    g0621(.A(new_n789), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G77), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n816), .A2(KEYINPUT32), .B1(G107), .B2(new_n810), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n818), .A2(new_n820), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n777), .B(new_n786), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n695), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n775), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n697), .A2(new_n786), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n695), .A2(G330), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  OAI22_X1  g0635(.A1(new_n789), .A2(new_n619), .B1(new_n798), .B2(new_n790), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n312), .B(new_n836), .C1(G294), .C2(new_n793), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G303), .A2(new_n802), .B1(new_n807), .B2(G107), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n809), .A2(new_n707), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n804), .B2(G283), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n820), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n809), .A2(new_n203), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n266), .B(new_n842), .C1(G132), .C2(new_n799), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n807), .A2(G50), .B1(new_n812), .B2(G58), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n793), .A2(G143), .B1(G159), .B2(new_n822), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(new_n804), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n801), .C1(new_n284), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n843), .B(new_n844), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n772), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n772), .A2(new_n773), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n785), .B1(new_n854), .B2(new_n215), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n347), .A2(new_n692), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n350), .B2(new_n351), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n346), .B1(new_n325), .B2(new_n326), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n329), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n329), .A3(new_n691), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n853), .B(new_n855), .C1(new_n863), .C2(new_n774), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n348), .A2(new_n352), .A3(new_n692), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n674), .A2(new_n675), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n751), .A2(new_n510), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n741), .B2(new_n862), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n739), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n785), .B1(new_n870), .B2(new_n739), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT103), .Z(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G384));
  INV_X1    g0675(.A(new_n553), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n876), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n230), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  NAND4_X1  g0680(.A1(new_n713), .A2(G77), .A3(new_n413), .A4(new_n414), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n277), .B(G13), .C1(new_n881), .C2(new_n250), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n425), .A2(new_n444), .ZN(new_n885));
  INV_X1    g0685(.A(new_n449), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n688), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n445), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT104), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n686), .B(KEYINPUT92), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n445), .B1(new_n459), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n893), .B2(new_n450), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n893), .C2(new_n450), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT79), .B1(new_n452), .B2(new_n453), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n460), .A2(new_n455), .A3(new_n461), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n888), .B1(new_n900), .B2(new_n446), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n884), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n892), .B1(new_n425), .B2(new_n444), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n463), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n895), .A2(new_n896), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(KEYINPUT38), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n377), .A2(new_n399), .A3(new_n691), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n658), .A2(new_n659), .A3(new_n446), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n903), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n888), .A2(KEYINPUT90), .A3(new_n445), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n425), .A2(new_n442), .A3(new_n444), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n903), .ZN(new_n914));
  AOI22_X1  g0714(.A1(KEYINPUT37), .A2(new_n912), .B1(new_n914), .B2(new_n887), .ZN(new_n915));
  NOR4_X1   g0715(.A1(new_n893), .A2(KEYINPUT90), .A3(new_n889), .A4(new_n450), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n463), .A2(new_n903), .B1(new_n895), .B2(new_n896), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(KEYINPUT38), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n907), .B(new_n909), .C1(new_n920), .C2(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n902), .A2(new_n906), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n399), .A2(new_n692), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n400), .A2(new_n403), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n403), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n399), .B(new_n692), .C1(new_n925), .C2(new_n377), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n868), .B2(new_n861), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n922), .A2(new_n929), .B1(new_n660), .B2(new_n892), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n464), .B1(new_n740), .B2(KEYINPUT29), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT105), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT105), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n743), .A2(new_n760), .A3(new_n936), .A4(new_n464), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n935), .A2(new_n667), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n932), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n736), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n730), .A2(new_n731), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n862), .B1(new_n926), .B2(new_n924), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT31), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n735), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT40), .B1(new_n920), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n922), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n464), .A3(new_n944), .A4(new_n941), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n911), .A2(new_n917), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n906), .B1(new_n952), .B2(KEYINPUT38), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n947), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT40), .B1(new_n902), .B2(new_n906), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(KEYINPUT40), .B1(new_n955), .B2(new_n947), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n941), .A2(new_n944), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n668), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n958), .A3(G330), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n939), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n277), .B2(new_n779), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n939), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n883), .B1(new_n961), .B2(new_n962), .ZN(G367));
  OAI211_X1 g0763(.A(new_n561), .B(new_n565), .C1(new_n559), .C2(new_n691), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n671), .A2(new_n692), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n702), .A2(new_n704), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n565), .B1(new_n964), .B2(new_n643), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n967), .A2(KEYINPUT42), .B1(new_n691), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n515), .A2(new_n691), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n517), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n669), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n968), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n966), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n703), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n711), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n702), .B(new_n704), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n984), .B2(new_n697), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(KEYINPUT107), .A3(new_n696), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(KEYINPUT108), .A3(new_n697), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n983), .B2(new_n696), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n761), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n705), .A2(new_n966), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT45), .Z(new_n994));
  NOR2_X1   g0794(.A1(new_n705), .A2(new_n966), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n996), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n994), .A2(new_n703), .A3(new_n996), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n703), .B1(new_n994), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n992), .B(new_n997), .C1(new_n1000), .C2(KEYINPUT106), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n981), .B1(new_n1001), .B2(new_n761), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n783), .ZN(new_n1003));
  INV_X1    g0803(.A(G143), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n801), .A2(new_n1004), .B1(new_n809), .B2(new_n215), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n312), .B1(new_n798), .B2(new_n846), .C1(new_n794), .C2(new_n284), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G58), .C2(new_n807), .ZN(new_n1007));
  INV_X1    g0807(.A(G159), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n847), .A2(new_n1008), .B1(new_n789), .B2(new_n201), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT109), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n819), .A2(G68), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n802), .A2(G311), .B1(G107), .B2(new_n812), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n206), .B2(new_n809), .C1(new_n592), .C2(new_n847), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n793), .A2(G303), .B1(G317), .B2(new_n799), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT46), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n806), .B2(new_n619), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n312), .B1(new_n822), .B2(G283), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1014), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n772), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n972), .A2(new_n775), .A3(new_n973), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n239), .A2(new_n765), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n776), .B(new_n1027), .C1(new_n211), .C2(new_n500), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n786), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1003), .A2(new_n1029), .ZN(G387));
  AOI22_X1  g0830(.A1(new_n709), .A2(new_n763), .B1(new_n207), .B2(new_n710), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n765), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G45), .B(new_n709), .C1(G68), .C2(G77), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n334), .A2(new_n201), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1038), .A2(KEYINPUT110), .B1(new_n244), .B2(new_n272), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1031), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n785), .B1(new_n1041), .B2(new_n776), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n775), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n702), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n806), .A2(new_n215), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n801), .A2(new_n1008), .B1(new_n809), .B2(new_n206), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n334), .C2(new_n804), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n819), .A2(new_n332), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n266), .B1(new_n799), .B2(G150), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n793), .A2(G50), .B1(G68), .B2(new_n822), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n312), .B1(new_n799), .B2(G326), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n793), .A2(G317), .B1(G303), .B2(new_n822), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n790), .B2(new_n847), .C1(new_n795), .C2(new_n801), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n807), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT49), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1052), .B1(new_n619), .B2(new_n809), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1060), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT111), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1051), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1044), .B1(new_n1065), .B2(new_n772), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n990), .B2(new_n783), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n991), .A2(new_n711), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n990), .A2(new_n761), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  OAI211_X1 g0870(.A(new_n1001), .B(new_n711), .C1(new_n992), .C2(new_n1000), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n978), .A2(new_n775), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n776), .B1(new_n206), .B2(new_n211), .C1(new_n248), .C2(new_n1032), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n786), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n794), .A2(new_n1008), .B1(new_n801), .B2(new_n284), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n819), .A2(G77), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n312), .B1(new_n798), .B2(new_n1004), .C1(new_n287), .C2(new_n789), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n839), .B1(new_n804), .B2(G50), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n203), .C2(new_n806), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n793), .A2(G311), .B1(new_n802), .B2(G317), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n804), .A2(G303), .B1(G107), .B2(new_n810), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n266), .B1(new_n798), .B2(new_n795), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G294), .B2(new_n822), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n807), .A2(G283), .B1(new_n812), .B2(G116), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1080), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n772), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1000), .A2(new_n783), .B1(new_n1072), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1071), .A2(new_n1094), .ZN(G390));
  OAI21_X1  g0895(.A(new_n907), .B1(new_n920), .B2(KEYINPUT39), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n773), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n785), .B1(new_n854), .B2(new_n287), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n789), .A2(new_n206), .B1(new_n798), .B2(new_n592), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n312), .B(new_n1099), .C1(G116), .C2(new_n793), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n847), .A2(new_n207), .B1(new_n538), .B2(new_n801), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1101), .A2(new_n815), .A3(new_n842), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n806), .A2(new_n284), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT53), .Z(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G159), .B2(new_n819), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n847), .A2(new_n846), .B1(new_n1107), .B2(new_n801), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n793), .A2(G132), .B1(G125), .B2(new_n799), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n266), .B1(new_n822), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1108), .B(new_n1113), .C1(G50), .C2(new_n810), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1103), .A2(new_n1079), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1097), .B(new_n1098), .C1(new_n827), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT114), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n929), .B2(new_n909), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n677), .A2(new_n865), .B1(new_n348), .B2(new_n691), .ZN(new_n1119));
  OAI211_X1 g0919(.A(KEYINPUT114), .B(new_n908), .C1(new_n1119), .C2(new_n928), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1096), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n908), .B(KEYINPUT113), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n920), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n759), .A2(new_n691), .A3(new_n860), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1124), .A2(new_n861), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n928), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n941), .A2(new_n942), .A3(G330), .A4(new_n944), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n732), .A2(new_n737), .A3(new_n863), .A4(new_n927), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1121), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1116), .B1(new_n1133), .B2(new_n780), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n941), .A2(G330), .A3(new_n944), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n928), .B1(new_n1135), .B2(new_n862), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1124), .A2(new_n1131), .A3(new_n861), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n732), .A2(new_n737), .A3(new_n863), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n928), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1128), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1119), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1136), .A2(new_n1137), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1135), .A2(new_n668), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n935), .A2(new_n937), .A3(new_n667), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n778), .B1(new_n1133), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1130), .A2(new_n1132), .A3(new_n1145), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1134), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(KEYINPUT118), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1144), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n302), .A2(new_n892), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n310), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n310), .A2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1154), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n1157), .A3(new_n1153), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n950), .B2(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n733), .B(new_n1165), .C1(new_n946), .C2(new_n949), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n931), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n956), .B2(new_n733), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n950), .A2(G330), .A3(new_n1163), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n932), .A3(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1148), .A2(new_n1152), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1151), .B1(new_n1171), .B2(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n778), .B1(new_n1171), .B2(KEYINPUT57), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1121), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1128), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1144), .B1(new_n1177), .B2(new_n1145), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1164), .A2(new_n1166), .A3(new_n931), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n932), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(KEYINPUT118), .B(new_n1174), .C1(new_n1178), .C2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1172), .A2(new_n1173), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1165), .A2(new_n773), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n312), .A2(G41), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1186), .B1(new_n538), .B2(new_n798), .C1(new_n794), .C2(new_n207), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n332), .B2(new_n822), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1045), .B1(G58), .B2(new_n810), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n804), .A2(G97), .B1(new_n802), .B2(G116), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n1012), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n793), .A2(G128), .B1(new_n807), .B2(new_n1111), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT115), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n819), .A2(G150), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n804), .A2(G132), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n802), .A2(G125), .B1(new_n822), .B2(G137), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT116), .Z(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1008), .B2(new_n809), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1203), .B2(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1196), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n827), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT117), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n785), .B(new_n1210), .C1(new_n201), .C2(new_n854), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1184), .A2(new_n783), .B1(new_n1185), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1183), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT119), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(G375));
  AND2_X1   g1015(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1216), .A2(new_n1145), .A3(new_n981), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n809), .A2(new_n215), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n801), .A2(new_n592), .B1(new_n806), .B2(new_n206), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G116), .C2(new_n804), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n312), .B1(new_n799), .B2(G303), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n793), .A2(G283), .B1(G107), .B2(new_n822), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n1048), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n789), .A2(new_n284), .B1(new_n798), .B2(new_n1107), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n266), .B(new_n1224), .C1(G137), .C2(new_n793), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n819), .A2(G50), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n802), .B1(new_n810), .B2(G58), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n804), .A2(new_n1111), .B1(G159), .B2(new_n807), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n827), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n785), .B(new_n1230), .C1(new_n203), .C2(new_n854), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n927), .B2(new_n774), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1142), .B2(new_n780), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1217), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G381));
  OR4_X1    g1035(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1236), .A2(G387), .A3(G381), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1214), .A3(new_n1149), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n689), .A2(G213), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT120), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(new_n1149), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT121), .ZN(G409));
  XNOR2_X1  g1044(.A(G393), .B(new_n834), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G387), .A2(new_n1247), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1246), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1239), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n711), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1142), .A2(new_n1144), .A3(KEYINPUT60), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT122), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1258), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1233), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G384), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n874), .A3(new_n1264), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1183), .A2(G378), .A3(new_n1212), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1171), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1212), .B1(new_n1271), .B2(new_n981), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1149), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1255), .B(new_n1269), .C1(new_n1270), .C2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1241), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(KEYINPUT126), .A3(new_n1241), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1275), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1240), .A2(G2897), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1266), .A2(new_n1267), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G2897), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1239), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT125), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1268), .A2(new_n1287), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1266), .B(new_n1267), .C1(new_n1286), .C2(new_n1241), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1279), .A2(new_n1280), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1254), .B1(new_n1283), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1276), .A2(new_n1239), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1295), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT123), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1274), .B2(KEYINPUT63), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OAI211_X1 g1107(.A(KEYINPUT123), .B(new_n1307), .C1(new_n1301), .C2(new_n1269), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1254), .A2(KEYINPUT61), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1300), .A2(new_n1304), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1299), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1213), .A2(G378), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1242), .A2(new_n1268), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1268), .B1(new_n1242), .B2(new_n1313), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1254), .B(KEYINPUT127), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1242), .A2(new_n1313), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1269), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1242), .A2(new_n1268), .A3(new_n1313), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1251), .A2(new_n1253), .A3(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1316), .A2(new_n1323), .ZN(G402));
endmodule


