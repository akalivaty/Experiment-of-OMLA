//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT11), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OR3_X1    g013(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT88), .A3(new_n211), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(G43gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(G50gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(G29gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT87), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G29gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(G36gat), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n223), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n216), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n223), .A2(new_n226), .A3(new_n231), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT89), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(KEYINPUT86), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(new_n211), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n226), .B1(new_n242), .B2(new_n231), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n209), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT90), .B(new_n243), .C1(new_n234), .C2(new_n237), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n208), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G15gat), .B(G22gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT16), .ZN(new_n249));
  AOI21_X1  g048(.A(G1gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G8gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n251), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT17), .A3(new_n244), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n252), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n251), .B(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n245), .B2(new_n246), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT18), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n256), .A2(KEYINPUT18), .A3(new_n257), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n233), .B1(new_n217), .B2(new_n232), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT89), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n244), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT90), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n238), .A2(new_n209), .A3(new_n244), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n254), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT13), .Z(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(KEYINPUT92), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT92), .B1(new_n272), .B2(new_n273), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n207), .B1(new_n265), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT92), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n207), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n264), .A4(new_n263), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n278), .A2(KEYINPUT93), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT93), .B1(new_n278), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G78gat), .B(G106gat), .Z(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT73), .B(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G148gat), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  OR3_X1    g091(.A1(new_n292), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n292), .B2(G148gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n300), .B2(KEYINPUT2), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n291), .A2(new_n302), .A3(new_n293), .A4(new_n294), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n296), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n297), .B(new_n300), .C1(new_n306), .C2(KEYINPUT2), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n304), .A2(new_n310), .A3(new_n305), .A4(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G211gat), .A2(G218gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(G211gat), .A2(G218gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n313), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT3), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n307), .B2(new_n304), .ZN(new_n326));
  OAI211_X1 g125(.A(G228gat), .B(G233gat), .C1(new_n323), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n321), .B(KEYINPUT78), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n307), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(KEYINPUT79), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n334), .B(new_n330), .C1(new_n329), .C2(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n336), .B(new_n337), .C1(new_n322), .C2(new_n312), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n327), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n327), .B2(new_n338), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n289), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT31), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n338), .A3(new_n339), .ZN(new_n345));
  INV_X1    g144(.A(new_n289), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n342), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n342), .B2(new_n347), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT24), .A3(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(KEYINPUT24), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT64), .ZN(new_n357));
  OR3_X1    g156(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT25), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT27), .B(G183gat), .Z(new_n363));
  OR3_X1    g162(.A1(new_n363), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT28), .B1(new_n363), .B2(G190gat), .ZN(new_n365));
  OR3_X1    g164(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(G176gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n366), .B(new_n367), .C1(new_n205), .C2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n364), .A2(new_n353), .A3(new_n365), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n356), .ZN(new_n371));
  NAND2_X1  g170(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n371), .B(new_n372), .C1(new_n360), .C2(KEYINPUT25), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n362), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT66), .B(G113gat), .Z(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT65), .B(G120gat), .ZN(new_n378));
  INV_X1    g177(.A(G113gat), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G127gat), .B(G134gat), .Z(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT1), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(G113gat), .B2(G120gat), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n380), .A2(new_n382), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n374), .A2(new_n385), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n390), .A3(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT32), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n389), .A2(new_n390), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G71gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n405), .B(G99gat), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n407), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n397), .A2(new_n400), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n351), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n374), .A2(new_n324), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT71), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n413), .A2(new_n415), .B1(new_n374), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n322), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n375), .A2(new_n415), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n374), .B2(new_n324), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n322), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424));
  INV_X1    g223(.A(G64gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G92gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n419), .A2(new_n422), .A3(new_n428), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n430), .A2(KEYINPUT72), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT72), .B1(new_n430), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT30), .B1(new_n423), .B2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n330), .A2(new_n386), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n304), .A2(new_n385), .A3(new_n307), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n309), .A2(new_n311), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n445), .A2(new_n386), .A3(new_n332), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(KEYINPUT4), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n304), .A2(new_n448), .A3(new_n385), .A4(new_n307), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n442), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n386), .A3(new_n332), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n453), .A2(new_n456), .A3(new_n438), .A4(new_n442), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT0), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G57gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G85gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n437), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n452), .B2(new_n457), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n437), .B(new_n464), .C1(new_n452), .C2(new_n457), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n434), .B(new_n436), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT35), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n342), .A2(new_n347), .ZN(new_n471));
  INV_X1    g270(.A(new_n348), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n342), .A2(new_n347), .A3(new_n348), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n436), .A2(new_n431), .A3(new_n430), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT84), .B1(new_n465), .B2(KEYINPUT6), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n462), .B(KEYINPUT80), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n458), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n452), .B2(new_n457), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n463), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n476), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n411), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n408), .A2(KEYINPUT85), .A3(new_n410), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n412), .A2(new_n470), .B1(new_n493), .B2(new_n469), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT83), .B(KEYINPUT38), .Z(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n423), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n428), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n423), .A2(new_n496), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n423), .A2(new_n429), .ZN(new_n501));
  OR3_X1    g300(.A1(new_n420), .A2(new_n421), .A3(new_n322), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(KEYINPUT37), .C1(new_n418), .C2(new_n417), .ZN(new_n503));
  INV_X1    g302(.A(new_n495), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n497), .A3(new_n428), .A4(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n480), .A2(new_n487), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n442), .B1(new_n453), .B2(new_n456), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT39), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n481), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n441), .A2(new_n443), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT81), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT40), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT81), .B(new_n517), .C1(new_n512), .C2(new_n514), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(new_n476), .A3(new_n485), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n475), .A2(new_n507), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT68), .B(KEYINPUT36), .Z(new_n521));
  AND3_X1   g320(.A1(new_n397), .A2(new_n400), .A3(new_n409), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n409), .B1(new_n397), .B2(new_n400), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT69), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n411), .A2(new_n526), .A3(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n408), .A2(KEYINPUT36), .A3(new_n410), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n408), .A2(KEYINPUT67), .A3(KEYINPUT36), .A4(new_n410), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n351), .A2(new_n468), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n288), .B1(new_n494), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(G85gat), .A3(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT8), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT98), .B(G92gat), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n542), .B(new_n544), .C1(G85gat), .C2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G92gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n427), .A2(KEYINPUT98), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(new_n547), .A3(new_n542), .A4(new_n544), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(KEYINPUT99), .A3(new_n548), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n557), .A2(KEYINPUT100), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT100), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n247), .A2(new_n255), .A3(new_n561), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n245), .A2(new_n246), .B1(new_n559), .B2(new_n560), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n562), .A2(new_n566), .A3(new_n563), .A4(new_n564), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(KEYINPUT97), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(KEYINPUT101), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n570), .A2(KEYINPUT101), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n577), .A3(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n573), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT21), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n425), .A2(G57gat), .ZN(new_n582));
  INV_X1    g381(.A(G57gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(G64gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT9), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  OR2_X1    g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n583), .B2(G64gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n425), .A2(KEYINPUT94), .A3(G57gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n590), .B1(new_n594), .B2(new_n582), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n254), .B1(new_n581), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT19), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n581), .ZN(new_n604));
  XOR2_X1   g403(.A(G183gat), .B(G211gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n603), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n580), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n556), .A2(new_n550), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n427), .A2(KEYINPUT98), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n552), .A2(G92gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n619), .A2(new_n551), .B1(KEYINPUT8), .B2(new_n543), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n547), .B1(new_n620), .B2(new_n542), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n558), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n557), .A2(KEYINPUT100), .A3(new_n558), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n614), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n557), .A2(new_n596), .A3(new_n558), .ZN(new_n627));
  INV_X1    g426(.A(new_n596), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n549), .A3(new_n556), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n627), .A2(new_n612), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n611), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n627), .A2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n611), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n368), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(G204gat), .Z(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n610), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n537), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n466), .A2(new_n467), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  INV_X1    g445(.A(G8gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n643), .B2(new_n476), .ZN(new_n648));
  INV_X1    g447(.A(new_n476), .ZN(new_n649));
  NOR2_X1   g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n249), .A2(new_n647), .ZN(new_n651));
  NOR4_X1   g450(.A1(new_n642), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n652), .ZN(G1325gat));
  AOI21_X1  g453(.A(G15gat), .B1(new_n643), .B2(new_n492), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT102), .Z(new_n656));
  INV_X1    g455(.A(new_n534), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n643), .A2(G15gat), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(G1326gat));
  OR3_X1    g458(.A1(new_n642), .A2(KEYINPUT103), .A3(new_n475), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT103), .B1(new_n642), .B2(new_n475), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT43), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(G22gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(G22gat), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n609), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n580), .A2(new_n640), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n537), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n228), .A2(new_n230), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n644), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(new_n644), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n493), .A2(new_n469), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n412), .A2(new_n470), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n536), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n580), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(KEYINPUT44), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n351), .B2(new_n468), .ZN(new_n684));
  AND4_X1   g483(.A1(KEYINPUT105), .A2(new_n473), .A3(new_n468), .A4(new_n474), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n520), .B(new_n534), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n580), .B1(new_n494), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n683), .B(new_n671), .C1(new_n687), .C2(KEYINPUT44), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n278), .A2(new_n284), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n640), .B(KEYINPUT104), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  INV_X1    g495(.A(new_n693), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n688), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n678), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n677), .B1(new_n700), .B2(new_n675), .ZN(G1328gat));
  NOR3_X1   g500(.A1(new_n673), .A2(G36gat), .A3(new_n649), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n649), .B1(new_n695), .B2(new_n699), .ZN(new_n704));
  INV_X1    g503(.A(G36gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(G1329gat));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n693), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n707), .B2(new_n534), .ZN(new_n708));
  INV_X1    g507(.A(new_n492), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n673), .A2(G43gat), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n657), .B1(new_n694), .B2(new_n698), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n707), .B2(new_n475), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n674), .A2(new_n221), .A3(new_n351), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n717), .ZN(new_n718));
  OR4_X1    g517(.A1(KEYINPUT107), .A2(new_n673), .A3(G50gat), .A4(new_n475), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n351), .B1(new_n694), .B2(new_n698), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G50gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n723), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g523(.A1(new_n494), .A2(new_n686), .ZN(new_n725));
  INV_X1    g524(.A(new_n692), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n610), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n691), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT108), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n678), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n583), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n729), .A2(new_n649), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  AND2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n732), .B2(new_n733), .ZN(G1333gat));
  NAND2_X1  g535(.A1(new_n657), .A2(G71gat), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n729), .A2(new_n709), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(G71gat), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT50), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n738), .B(new_n742), .C1(G71gat), .C2(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n475), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT109), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  OR2_X1    g546(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n609), .A2(new_n690), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n640), .A3(new_n683), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n678), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n725), .A2(new_n682), .A3(new_n749), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n687), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n756), .A2(G85gat), .A3(new_n678), .ZN(new_n757));
  INV_X1    g556(.A(new_n640), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  OAI21_X1  g558(.A(new_n545), .B1(new_n750), .B2(new_n649), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n726), .A2(G92gat), .A3(new_n649), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n760), .B(new_n761), .C1(new_n756), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n754), .A2(new_n765), .A3(new_n755), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n753), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n762), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n767), .A4(new_n762), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n770), .A2(new_n760), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n764), .B1(new_n772), .B2(new_n761), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n750), .B2(new_n534), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n756), .A2(G99gat), .A3(new_n709), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n758), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n475), .A2(G106gat), .A3(new_n726), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(G106gat), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n683), .B(new_n749), .C1(new_n687), .C2(KEYINPUT44), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(new_n475), .A3(new_n758), .ZN(new_n782));
  OAI221_X1 g581(.A(new_n777), .B1(new_n756), .B2(new_n779), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT112), .B(G106gat), .C1(new_n750), .C2(new_n475), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n782), .B2(new_n780), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n767), .A3(new_n778), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n788), .B2(new_n777), .ZN(G1339gat));
  AND4_X1   g588(.A1(new_n691), .A2(new_n580), .A3(new_n609), .A4(new_n758), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n613), .B1(new_n559), .B2(new_n560), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n627), .A2(new_n612), .A3(new_n629), .ZN(new_n792));
  INV_X1    g591(.A(new_n611), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n631), .A2(new_n794), .A3(KEYINPUT113), .A4(KEYINPUT54), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n636), .B1(new_n631), .B2(KEYINPUT54), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(new_n800), .C1(new_n797), .C2(new_n798), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n804), .A3(new_n637), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n570), .A2(KEYINPUT101), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n578), .A3(new_n573), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n257), .B1(new_n256), .B2(new_n260), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n272), .A2(new_n273), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n206), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n284), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n805), .A2(new_n807), .A3(new_n575), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n284), .A2(new_n640), .A3(new_n810), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n805), .B2(new_n690), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n682), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT114), .B(new_n790), .C1(new_n815), .C2(new_n671), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n804), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n690), .A2(new_n818), .A3(new_n638), .ZN(new_n819));
  INV_X1    g618(.A(new_n813), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n819), .A2(new_n820), .B1(new_n807), .B2(new_n575), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n801), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n803), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n638), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n284), .A2(new_n810), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n580), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n671), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n790), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n817), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n709), .A2(new_n351), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n678), .A2(new_n476), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n288), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT115), .Z(new_n836));
  AND3_X1   g635(.A1(new_n831), .A2(new_n412), .A3(new_n833), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n691), .A2(new_n376), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT116), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n834), .B2(new_n726), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(new_n378), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n837), .A2(new_n844), .A3(new_n640), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n834), .A2(new_n847), .A3(new_n671), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT118), .Z(new_n849));
  AOI21_X1  g648(.A(G127gat), .B1(new_n837), .B2(new_n609), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n852), .A3(new_n682), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT56), .Z(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n834), .B2(new_n580), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n534), .A2(new_n833), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n831), .A2(new_n351), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(G141gat), .A3(new_n288), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n475), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n285), .A2(new_n286), .A3(new_n825), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n580), .B1(new_n865), .B2(new_n813), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n609), .B1(new_n866), .B2(new_n812), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n867), .B2(new_n790), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n864), .C1(new_n867), .C2(new_n790), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n828), .A2(new_n829), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT114), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n828), .A2(new_n817), .A3(new_n829), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n863), .B1(new_n876), .B2(new_n475), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n858), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n287), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n857), .B(new_n862), .C1(new_n879), .C2(new_n290), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n869), .A2(new_n871), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n831), .B2(new_n351), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n690), .B(new_n859), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n290), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n862), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n887), .B2(KEYINPUT58), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n861), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT120), .A3(new_n857), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n880), .B1(new_n888), .B2(new_n890), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n475), .ZN(new_n892));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n858), .A2(new_n758), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n640), .B(new_n859), .C1(new_n882), .C2(new_n883), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(G148gat), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n896), .A2(KEYINPUT121), .A3(new_n897), .A4(G148gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n875), .A3(new_n864), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT122), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n831), .A2(new_n905), .A3(new_n864), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n287), .A2(new_n610), .A3(new_n640), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n351), .B1(new_n867), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n863), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n894), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n893), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n894), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n897), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n895), .B1(new_n902), .B2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(new_n298), .B1(new_n878), .B2(new_n609), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n860), .A2(G155gat), .A3(new_n671), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  NAND4_X1  g721(.A1(new_n892), .A2(new_n299), .A3(new_n682), .A4(new_n859), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n878), .A2(new_n682), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n299), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n644), .A2(new_n649), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n876), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n832), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n288), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n412), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n690), .A2(new_n205), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  NOR3_X1   g732(.A1(new_n929), .A2(new_n368), .A3(new_n726), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n412), .A3(new_n640), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n368), .B2(new_n935), .ZN(G1349gat));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n929), .B2(new_n671), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n671), .A2(new_n363), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n928), .A2(new_n412), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(KEYINPUT60), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n929), .B2(new_n580), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n580), .A2(G190gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n931), .B2(new_n951), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n910), .A2(new_n534), .A3(new_n926), .ZN(new_n953));
  OAI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n288), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n657), .A2(new_n927), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n892), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n690), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n892), .A2(new_n958), .A3(new_n955), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT126), .B1(new_n960), .B2(new_n691), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n954), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n892), .A2(new_n955), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(G204gat), .A3(new_n758), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n953), .B2(new_n726), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1353gat));
  OR3_X1    g771(.A1(new_n968), .A2(G211gat), .A3(new_n671), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n910), .A2(new_n534), .A3(new_n609), .A4(new_n926), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n953), .A2(new_n978), .A3(new_n580), .ZN(new_n979));
  AOI21_X1  g778(.A(G218gat), .B1(new_n956), .B2(new_n682), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(G1355gat));
endmodule


