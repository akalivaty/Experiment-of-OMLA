

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776;

  AND2_X1 U372 ( .A1(n388), .A2(n662), .ZN(n358) );
  AND2_X1 U373 ( .A1(n654), .A2(G472), .ZN(n360) );
  NOR2_X1 U374 ( .A1(n636), .A2(n613), .ZN(n681) );
  INV_X1 U375 ( .A(n430), .ZN(n351) );
  INV_X1 U376 ( .A(KEYINPUT88), .ZN(n350) );
  BUF_X1 U377 ( .A(G107), .Z(n676) );
  INV_X2 U378 ( .A(n397), .ZN(n390) );
  XNOR2_X2 U379 ( .A(n404), .B(KEYINPUT83), .ZN(n764) );
  XNOR2_X2 U380 ( .A(n559), .B(KEYINPUT105), .ZN(n619) );
  XNOR2_X2 U381 ( .A(n475), .B(n474), .ZN(n745) );
  NAND2_X1 U382 ( .A1(n351), .A2(n350), .ZN(n352) );
  AND2_X2 U383 ( .A1(n423), .A2(n352), .ZN(n420) );
  NOR2_X4 U384 ( .A1(n688), .A2(n653), .ZN(n691) );
  INV_X2 U385 ( .A(G953), .ZN(n765) );
  OR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n354) );
  NOR2_X2 U387 ( .A1(n742), .A2(n749), .ZN(n743) );
  AND2_X2 U388 ( .A1(n377), .A2(n376), .ZN(n381) );
  INV_X1 U389 ( .A(n539), .ZN(n562) );
  AND2_X1 U390 ( .A1(n386), .A2(n389), .ZN(n385) );
  NAND2_X1 U391 ( .A1(n405), .A2(n366), .ZN(n404) );
  NOR2_X1 U392 ( .A1(n626), .A2(n625), .ZN(n638) );
  NAND2_X1 U393 ( .A1(n420), .A2(n417), .ZN(n530) );
  AND2_X1 U394 ( .A1(n704), .A2(n703), .ZN(n591) );
  BUF_X1 U395 ( .A(n559), .Z(n701) );
  XNOR2_X1 U396 ( .A(n441), .B(n440), .ZN(n559) );
  XNOR2_X1 U397 ( .A(n739), .B(n738), .ZN(n740) );
  OR2_X1 U398 ( .A1(n664), .A2(G902), .ZN(n525) );
  XNOR2_X1 U399 ( .A(n415), .B(n414), .ZN(n539) );
  XNOR2_X1 U400 ( .A(n454), .B(n455), .ZN(n747) );
  XNOR2_X1 U401 ( .A(KEYINPUT16), .B(G122), .ZN(n498) );
  INV_X1 U402 ( .A(G210), .ZN(n363) );
  NAND2_X1 U403 ( .A1(n397), .A2(n357), .ZN(n355) );
  AND2_X1 U404 ( .A1(n355), .A2(n356), .ZN(n386) );
  OR2_X1 U405 ( .A1(n662), .A2(n391), .ZN(n356) );
  AND2_X1 U406 ( .A1(n372), .A2(n394), .ZN(n357) );
  AND2_X4 U407 ( .A1(n408), .A2(n654), .ZN(n397) );
  AND2_X1 U408 ( .A1(n395), .A2(n364), .ZN(G63) );
  XNOR2_X1 U409 ( .A(n745), .B(n744), .ZN(n364) );
  AND2_X1 U410 ( .A1(n393), .A2(n391), .ZN(n359) );
  NAND2_X1 U411 ( .A1(n408), .A2(n360), .ZN(n384) );
  BUF_X1 U412 ( .A(n602), .Z(n361) );
  XNOR2_X1 U413 ( .A(n549), .B(KEYINPUT35), .ZN(n602) );
  NAND2_X1 U414 ( .A1(n408), .A2(n362), .ZN(n741) );
  NOR2_X1 U415 ( .A1(n691), .A2(n363), .ZN(n362) );
  XNOR2_X2 U416 ( .A(n399), .B(n756), .ZN(n736) );
  AND2_X1 U417 ( .A1(n430), .A2(KEYINPUT88), .ZN(n418) );
  NOR2_X1 U418 ( .A1(n426), .A2(n716), .ZN(n425) );
  XNOR2_X1 U419 ( .A(n643), .B(KEYINPUT46), .ZN(n412) );
  XNOR2_X1 U420 ( .A(n470), .B(n479), .ZN(n516) );
  NAND2_X1 U421 ( .A1(n765), .A2(G224), .ZN(n500) );
  XNOR2_X1 U422 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n621) );
  INV_X1 U423 ( .A(KEYINPUT110), .ZN(n617) );
  OR2_X1 U424 ( .A1(n511), .A2(n650), .ZN(n428) );
  XOR2_X1 U425 ( .A(KEYINPUT98), .B(KEYINPUT81), .Z(n446) );
  XNOR2_X1 U426 ( .A(G128), .B(G119), .ZN(n444) );
  XNOR2_X1 U427 ( .A(G140), .B(KEYINPUT10), .ZN(n448) );
  XNOR2_X1 U428 ( .A(n450), .B(n411), .ZN(n410) );
  INV_X1 U429 ( .A(KEYINPUT8), .ZN(n411) );
  NAND2_X1 U430 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  XNOR2_X1 U431 ( .A(n407), .B(n604), .ZN(n406) );
  INV_X1 U432 ( .A(n404), .ZN(n652) );
  XNOR2_X1 U433 ( .A(n456), .B(n365), .ZN(n414) );
  OR2_X1 U434 ( .A1(n747), .A2(G902), .ZN(n415) );
  XNOR2_X1 U435 ( .A(G113), .B(G122), .ZN(n482) );
  XNOR2_X1 U436 ( .A(G104), .B(G143), .ZN(n483) );
  XNOR2_X1 U437 ( .A(KEYINPUT68), .B(G131), .ZN(n479) );
  XNOR2_X1 U438 ( .A(G137), .B(KEYINPUT5), .ZN(n432) );
  XOR2_X1 U439 ( .A(KEYINPUT24), .B(G110), .Z(n445) );
  INV_X1 U440 ( .A(G134), .ZN(n431) );
  XNOR2_X1 U441 ( .A(KEYINPUT69), .B(G137), .ZN(n515) );
  NAND2_X1 U442 ( .A1(n750), .A2(n650), .ZN(n407) );
  INV_X1 U443 ( .A(KEYINPUT82), .ZN(n604) );
  XNOR2_X1 U444 ( .A(n646), .B(n370), .ZN(n405) );
  INV_X1 U445 ( .A(G237), .ZN(n508) );
  NAND2_X1 U446 ( .A1(n511), .A2(n650), .ZN(n429) );
  XNOR2_X1 U447 ( .A(G116), .B(G122), .ZN(n468) );
  XNOR2_X1 U448 ( .A(n501), .B(n502), .ZN(n403) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n458) );
  NAND2_X1 U450 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U451 ( .A(n618), .B(n617), .ZN(n624) );
  XNOR2_X1 U452 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U453 ( .A(n449), .B(n761), .ZN(n455) );
  NOR2_X1 U454 ( .A1(n392), .A2(n749), .ZN(n391) );
  NOR2_X1 U455 ( .A1(n396), .A2(G475), .ZN(n392) );
  BUF_X1 U456 ( .A(G101), .Z(n398) );
  XOR2_X1 U457 ( .A(n457), .B(KEYINPUT79), .Z(n365) );
  AND2_X1 U458 ( .A1(n775), .A2(n649), .ZN(n366) );
  AND2_X1 U459 ( .A1(n578), .A2(n577), .ZN(n367) );
  NOR2_X1 U460 ( .A1(n773), .A2(KEYINPUT44), .ZN(n368) );
  AND2_X1 U461 ( .A1(n427), .A2(n429), .ZN(n369) );
  XOR2_X1 U462 ( .A(KEYINPUT48), .B(KEYINPUT84), .Z(n370) );
  INV_X1 U463 ( .A(n661), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U465 ( .A(KEYINPUT62), .B(n655), .ZN(n371) );
  AND2_X1 U466 ( .A1(n396), .A2(G475), .ZN(n372) );
  AND2_X1 U467 ( .A1(n661), .A2(n394), .ZN(n373) );
  XNOR2_X1 U468 ( .A(n657), .B(KEYINPUT89), .ZN(n374) );
  XOR2_X1 U469 ( .A(G110), .B(KEYINPUT117), .Z(n375) );
  AND2_X1 U470 ( .A1(n656), .A2(G953), .ZN(n749) );
  INV_X1 U471 ( .A(n749), .ZN(n395) );
  INV_X1 U472 ( .A(n662), .ZN(n394) );
  AND2_X1 U473 ( .A1(n668), .A2(n599), .ZN(n376) );
  NAND2_X1 U474 ( .A1(n582), .A2(n581), .ZN(n377) );
  XNOR2_X2 U475 ( .A(n378), .B(KEYINPUT45), .ZN(n750) );
  NAND2_X1 U476 ( .A1(n381), .A2(n379), .ZN(n378) );
  NAND2_X1 U477 ( .A1(n380), .A2(n603), .ZN(n379) );
  NAND2_X1 U478 ( .A1(n601), .A2(n600), .ZN(n380) );
  XNOR2_X1 U479 ( .A(n382), .B(n374), .ZN(G57) );
  NAND2_X1 U480 ( .A1(n383), .A2(n395), .ZN(n382) );
  XNOR2_X1 U481 ( .A(n384), .B(n371), .ZN(n383) );
  NAND2_X1 U482 ( .A1(n387), .A2(n385), .ZN(G60) );
  NAND2_X1 U483 ( .A1(n358), .A2(n359), .ZN(n387) );
  NAND2_X1 U484 ( .A1(n397), .A2(n372), .ZN(n393) );
  NAND2_X1 U485 ( .A1(n390), .A2(n661), .ZN(n388) );
  NAND2_X1 U486 ( .A1(n390), .A2(n373), .ZN(n389) );
  XNOR2_X1 U487 ( .A(n530), .B(n529), .ZN(n612) );
  NAND2_X1 U488 ( .A1(n572), .A2(n556), .ZN(n558) );
  XNOR2_X1 U489 ( .A(n555), .B(n554), .ZN(n572) );
  XNOR2_X2 U490 ( .A(n517), .B(n498), .ZN(n401) );
  XNOR2_X1 U491 ( .A(n400), .B(n403), .ZN(n399) );
  XNOR2_X1 U492 ( .A(n402), .B(n506), .ZN(n400) );
  XNOR2_X2 U493 ( .A(n401), .B(n499), .ZN(n756) );
  XNOR2_X1 U494 ( .A(n500), .B(n503), .ZN(n402) );
  XNOR2_X2 U495 ( .A(n497), .B(G104), .ZN(n517) );
  NAND2_X1 U496 ( .A1(n406), .A2(n764), .ZN(n409) );
  INV_X1 U497 ( .A(n750), .ZN(n688) );
  NAND2_X2 U498 ( .A1(n409), .A2(n651), .ZN(n408) );
  NAND2_X1 U499 ( .A1(n424), .A2(n513), .ZN(n423) );
  XNOR2_X2 U500 ( .A(n609), .B(n526), .ZN(n704) );
  NAND2_X1 U501 ( .A1(n410), .A2(G221), .ZN(n453) );
  NAND2_X1 U502 ( .A1(n410), .A2(G217), .ZN(n473) );
  NAND2_X1 U503 ( .A1(n413), .A2(n412), .ZN(n646) );
  AND2_X1 U504 ( .A1(n645), .A2(n644), .ZN(n413) );
  NAND2_X1 U505 ( .A1(n579), .A2(n368), .ZN(n601) );
  XNOR2_X1 U506 ( .A(n579), .B(n375), .ZN(G12) );
  XNOR2_X2 U507 ( .A(n564), .B(n416), .ZN(n579) );
  INV_X1 U508 ( .A(KEYINPUT107), .ZN(n416) );
  NAND2_X1 U509 ( .A1(n736), .A2(n511), .ZN(n430) );
  INV_X1 U510 ( .A(n424), .ZN(n419) );
  NAND2_X1 U511 ( .A1(n369), .A2(n430), .ZN(n568) );
  NAND2_X1 U512 ( .A1(n427), .A2(n425), .ZN(n424) );
  INV_X1 U513 ( .A(n429), .ZN(n426) );
  OR2_X2 U514 ( .A1(n736), .A2(n428), .ZN(n427) );
  NAND2_X1 U515 ( .A1(n591), .A2(n570), .ZN(n542) );
  INV_X1 U516 ( .A(KEYINPUT28), .ZN(n606) );
  XNOR2_X1 U517 ( .A(n606), .B(KEYINPUT113), .ZN(n607) );
  XNOR2_X1 U518 ( .A(n516), .B(n515), .ZN(n763) );
  XNOR2_X1 U519 ( .A(n608), .B(n607), .ZN(n611) );
  BUF_X1 U520 ( .A(n612), .Z(n613) );
  XNOR2_X2 U521 ( .A(G143), .B(G128), .ZN(n505) );
  XNOR2_X1 U522 ( .A(n505), .B(n431), .ZN(n470) );
  XNOR2_X2 U523 ( .A(KEYINPUT4), .B(G101), .ZN(n503) );
  XNOR2_X1 U524 ( .A(n503), .B(G146), .ZN(n522) );
  XNOR2_X1 U525 ( .A(n432), .B(KEYINPUT76), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n522), .B(n433), .ZN(n438) );
  XNOR2_X1 U527 ( .A(KEYINPUT77), .B(n354), .ZN(n478) );
  NAND2_X1 U528 ( .A1(n478), .A2(G210), .ZN(n436) );
  XNOR2_X1 U529 ( .A(G116), .B(G113), .ZN(n435) );
  XNOR2_X1 U530 ( .A(KEYINPUT3), .B(G119), .ZN(n434) );
  XNOR2_X1 U531 ( .A(n435), .B(n434), .ZN(n499) );
  XNOR2_X1 U532 ( .A(n436), .B(n499), .ZN(n437) );
  XNOR2_X1 U533 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U534 ( .A(n516), .B(n439), .ZN(n655) );
  INV_X1 U535 ( .A(G902), .ZN(n509) );
  NAND2_X1 U536 ( .A1(n655), .A2(n509), .ZN(n441) );
  XOR2_X1 U537 ( .A(G472), .B(KEYINPUT73), .Z(n440) );
  INV_X1 U538 ( .A(KEYINPUT6), .ZN(n442) );
  XNOR2_X1 U539 ( .A(n701), .B(n442), .ZN(n570) );
  XNOR2_X1 U540 ( .A(G902), .B(KEYINPUT15), .ZN(n507) );
  NAND2_X1 U541 ( .A1(n507), .A2(G234), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n443), .B(KEYINPUT20), .ZN(n463) );
  NAND2_X1 U543 ( .A1(n463), .A2(G217), .ZN(n456) );
  XNOR2_X1 U544 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U545 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X2 U546 ( .A(G146), .B(G125), .ZN(n504) );
  XNOR2_X1 U547 ( .A(n504), .B(n448), .ZN(n761) );
  NAND2_X1 U548 ( .A1(G234), .A2(n765), .ZN(n450) );
  INV_X1 U549 ( .A(n515), .ZN(n451) );
  XOR2_X1 U550 ( .A(n451), .B(KEYINPUT23), .Z(n452) );
  XNOR2_X1 U551 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n457) );
  XOR2_X1 U553 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n459) );
  XNOR2_X1 U554 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U555 ( .A1(G952), .A2(n460), .ZN(n732) );
  NOR2_X1 U556 ( .A1(n732), .A2(G953), .ZN(n534) );
  NAND2_X1 U557 ( .A1(G902), .A2(n460), .ZN(n532) );
  OR2_X1 U558 ( .A1(n765), .A2(n532), .ZN(n461) );
  NOR2_X1 U559 ( .A1(G900), .A2(n461), .ZN(n462) );
  NOR2_X1 U560 ( .A1(n534), .A2(n462), .ZN(n626) );
  AND2_X1 U561 ( .A1(n463), .A2(G221), .ZN(n464) );
  XNOR2_X1 U562 ( .A(n464), .B(KEYINPUT21), .ZN(n698) );
  INV_X1 U563 ( .A(n698), .ZN(n465) );
  NOR2_X1 U564 ( .A1(n626), .A2(n465), .ZN(n466) );
  NAND2_X1 U565 ( .A1(n562), .A2(n466), .ZN(n467) );
  XNOR2_X1 U566 ( .A(n467), .B(KEYINPUT70), .ZN(n605) );
  XNOR2_X1 U567 ( .A(n468), .B(n676), .ZN(n469) );
  XOR2_X1 U568 ( .A(n469), .B(KEYINPUT9), .Z(n472) );
  INV_X1 U569 ( .A(n470), .ZN(n471) );
  XNOR2_X1 U570 ( .A(n472), .B(n471), .ZN(n475) );
  XNOR2_X1 U571 ( .A(n473), .B(KEYINPUT7), .ZN(n474) );
  NAND2_X1 U572 ( .A1(n745), .A2(n509), .ZN(n477) );
  INV_X1 U573 ( .A(G478), .ZN(n476) );
  XNOR2_X1 U574 ( .A(n477), .B(n476), .ZN(n595) );
  NAND2_X1 U575 ( .A1(n478), .A2(G214), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U577 ( .A(n761), .B(n481), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U579 ( .A(KEYINPUT101), .B(KEYINPUT11), .ZN(n485) );
  XNOR2_X1 U580 ( .A(KEYINPUT12), .B(KEYINPUT100), .ZN(n484) );
  XNOR2_X1 U581 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U583 ( .A(n489), .B(n488), .ZN(n660) );
  OR2_X1 U584 ( .A1(n660), .A2(G902), .ZN(n492) );
  XNOR2_X1 U585 ( .A(KEYINPUT13), .B(G475), .ZN(n490) );
  XNOR2_X1 U586 ( .A(n490), .B(KEYINPUT102), .ZN(n491) );
  XNOR2_X1 U587 ( .A(n492), .B(n491), .ZN(n550) );
  INV_X1 U588 ( .A(n550), .ZN(n594) );
  NAND2_X1 U589 ( .A1(n595), .A2(n594), .ZN(n641) );
  INV_X1 U590 ( .A(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n641), .B(n493), .ZN(n683) );
  INV_X1 U592 ( .A(n683), .ZN(n494) );
  NOR2_X1 U593 ( .A1(n605), .A2(n494), .ZN(n495) );
  NAND2_X1 U594 ( .A1(n570), .A2(n495), .ZN(n496) );
  XNOR2_X1 U595 ( .A(KEYINPUT109), .B(n496), .ZN(n565) );
  XNOR2_X2 U596 ( .A(G110), .B(G107), .ZN(n497) );
  XNOR2_X1 U597 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n501) );
  XNOR2_X1 U598 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n502) );
  XNOR2_X1 U599 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U600 ( .A(n507), .ZN(n650) );
  NAND2_X1 U601 ( .A1(n509), .A2(n508), .ZN(n512) );
  NAND2_X1 U602 ( .A1(n512), .A2(G210), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n510), .B(KEYINPUT94), .ZN(n511) );
  NAND2_X1 U604 ( .A1(n512), .A2(G214), .ZN(n632) );
  INV_X1 U605 ( .A(n632), .ZN(n716) );
  INV_X1 U606 ( .A(KEYINPUT88), .ZN(n513) );
  NAND2_X1 U607 ( .A1(n565), .A2(n530), .ZN(n514) );
  XOR2_X1 U608 ( .A(KEYINPUT36), .B(n514), .Z(n527) );
  BUF_X1 U609 ( .A(n517), .Z(n518) );
  INV_X1 U610 ( .A(n518), .ZN(n521) );
  NAND2_X1 U611 ( .A1(n765), .A2(G227), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(G140), .ZN(n520) );
  XNOR2_X1 U613 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U614 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U615 ( .A(n763), .B(n524), .ZN(n664) );
  XNOR2_X2 U616 ( .A(n525), .B(G469), .ZN(n609) );
  XNOR2_X1 U617 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n526) );
  NAND2_X1 U618 ( .A1(n527), .A2(n704), .ZN(n644) );
  XOR2_X1 U619 ( .A(G125), .B(KEYINPUT37), .Z(n528) );
  XNOR2_X1 U620 ( .A(n644), .B(n528), .ZN(G27) );
  XNOR2_X1 U621 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n529) );
  NOR2_X1 U622 ( .A1(G898), .A2(n765), .ZN(n531) );
  XNOR2_X1 U623 ( .A(KEYINPUT95), .B(n531), .ZN(n757) );
  NOR2_X1 U624 ( .A1(n532), .A2(n757), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n533), .B(KEYINPUT96), .ZN(n535) );
  NOR2_X1 U626 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X2 U627 ( .A1(n612), .A2(n536), .ZN(n537) );
  XNOR2_X2 U628 ( .A(n537), .B(KEYINPUT0), .ZN(n590) );
  INV_X1 U629 ( .A(n590), .ZN(n538) );
  XNOR2_X1 U630 ( .A(n538), .B(KEYINPUT97), .ZN(n589) );
  AND2_X1 U631 ( .A1(n698), .A2(n539), .ZN(n703) );
  XNOR2_X1 U632 ( .A(KEYINPUT91), .B(KEYINPUT33), .ZN(n540) );
  XNOR2_X1 U633 ( .A(n540), .B(KEYINPUT71), .ZN(n541) );
  XNOR2_X1 U634 ( .A(n542), .B(n541), .ZN(n693) );
  NAND2_X1 U635 ( .A1(n589), .A2(n693), .ZN(n544) );
  XNOR2_X1 U636 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n543) );
  XNOR2_X1 U637 ( .A(n544), .B(n543), .ZN(n545) );
  INV_X1 U638 ( .A(n545), .ZN(n548) );
  INV_X1 U639 ( .A(n595), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n546), .A2(n594), .ZN(n627) );
  INV_X1 U641 ( .A(n627), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U643 ( .A(G122), .B(n361), .Z(G24) );
  NAND2_X1 U644 ( .A1(n595), .A2(n550), .ZN(n552) );
  INV_X1 U645 ( .A(KEYINPUT104), .ZN(n551) );
  XNOR2_X1 U646 ( .A(n552), .B(n551), .ZN(n718) );
  AND2_X1 U647 ( .A1(n718), .A2(n698), .ZN(n553) );
  NAND2_X1 U648 ( .A1(n590), .A2(n553), .ZN(n555) );
  INV_X1 U649 ( .A(KEYINPUT22), .ZN(n554) );
  INV_X1 U650 ( .A(n704), .ZN(n556) );
  INV_X1 U651 ( .A(KEYINPUT106), .ZN(n557) );
  XNOR2_X1 U652 ( .A(n558), .B(n557), .ZN(n560) );
  NAND2_X1 U653 ( .A1(n560), .A2(n619), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n561), .B(KEYINPUT65), .ZN(n563) );
  NAND2_X1 U655 ( .A1(n563), .A2(n562), .ZN(n564) );
  AND2_X1 U656 ( .A1(n565), .A2(n632), .ZN(n566) );
  NAND2_X1 U657 ( .A1(n566), .A2(n556), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n567), .B(KEYINPUT43), .ZN(n569) );
  NAND2_X1 U659 ( .A1(n569), .A2(n568), .ZN(n649) );
  XNOR2_X1 U660 ( .A(n649), .B(G140), .ZN(G42) );
  INV_X1 U661 ( .A(KEYINPUT87), .ZN(n600) );
  NAND2_X1 U662 ( .A1(n602), .A2(n600), .ZN(n578) );
  INV_X1 U663 ( .A(n570), .ZN(n571) );
  AND2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n583) );
  AND2_X1 U665 ( .A1(n704), .A2(n562), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n583), .A2(n573), .ZN(n576) );
  INV_X1 U667 ( .A(KEYINPUT64), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n574), .B(KEYINPUT32), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n576), .B(n575), .ZN(n773) );
  INV_X1 U670 ( .A(KEYINPUT44), .ZN(n580) );
  NOR2_X1 U671 ( .A1(n773), .A2(n580), .ZN(n577) );
  NAND2_X1 U672 ( .A1(n579), .A2(n367), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n600), .A2(n580), .ZN(n581) );
  XNOR2_X1 U674 ( .A(n583), .B(KEYINPUT85), .ZN(n584) );
  OR2_X1 U675 ( .A1(n584), .A2(n704), .ZN(n586) );
  INV_X1 U676 ( .A(KEYINPUT86), .ZN(n585) );
  XNOR2_X1 U677 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U678 ( .A1(n587), .A2(n539), .ZN(n668) );
  NAND2_X1 U679 ( .A1(n703), .A2(n609), .ZN(n618) );
  NOR2_X1 U680 ( .A1(n618), .A2(n701), .ZN(n588) );
  AND2_X1 U681 ( .A1(n589), .A2(n588), .ZN(n672) );
  BUF_X1 U682 ( .A(n590), .Z(n592) );
  AND2_X1 U683 ( .A1(n591), .A2(n701), .ZN(n709) );
  NAND2_X1 U684 ( .A1(n592), .A2(n709), .ZN(n593) );
  XNOR2_X1 U685 ( .A(n593), .B(KEYINPUT31), .ZN(n686) );
  OR2_X1 U686 ( .A1(n672), .A2(n686), .ZN(n596) );
  OR2_X1 U687 ( .A1(n595), .A2(n594), .ZN(n671) );
  AND2_X1 U688 ( .A1(n671), .A2(n641), .ZN(n722) );
  INV_X1 U689 ( .A(n722), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n596), .A2(n614), .ZN(n598) );
  INV_X1 U691 ( .A(KEYINPUT103), .ZN(n597) );
  XNOR2_X1 U692 ( .A(n598), .B(n597), .ZN(n599) );
  INV_X1 U693 ( .A(n361), .ZN(n603) );
  NOR2_X1 U694 ( .A1(n605), .A2(n619), .ZN(n608) );
  XNOR2_X1 U695 ( .A(n609), .B(KEYINPUT112), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n636) );
  NAND2_X1 U697 ( .A1(n681), .A2(n614), .ZN(n615) );
  NOR2_X1 U698 ( .A1(KEYINPUT67), .A2(n615), .ZN(n616) );
  XNOR2_X1 U699 ( .A(KEYINPUT47), .B(n616), .ZN(n629) );
  INV_X1 U700 ( .A(n619), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n620), .A2(n632), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n627), .A2(n568), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n638), .A2(n628), .ZN(n680) );
  NAND2_X1 U705 ( .A1(n629), .A2(n680), .ZN(n631) );
  INV_X1 U706 ( .A(KEYINPUT74), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n645) );
  XNOR2_X1 U708 ( .A(n568), .B(KEYINPUT38), .ZN(n715) );
  NAND2_X1 U709 ( .A1(n715), .A2(n632), .ZN(n721) );
  INV_X1 U710 ( .A(n721), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n633), .A2(n718), .ZN(n635) );
  INV_X1 U712 ( .A(KEYINPUT41), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n635), .B(n634), .ZN(n713) );
  NOR2_X1 U714 ( .A1(n636), .A2(n713), .ZN(n637) );
  XNOR2_X1 U715 ( .A(KEYINPUT42), .B(n637), .ZN(n776) );
  NAND2_X1 U716 ( .A1(n638), .A2(n715), .ZN(n640) );
  INV_X1 U717 ( .A(KEYINPUT39), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n640), .B(n639), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n647), .A2(n641), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT40), .ZN(n774) );
  NOR2_X1 U721 ( .A1(n776), .A2(n774), .ZN(n643) );
  OR2_X1 U722 ( .A1(n647), .A2(n671), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(KEYINPUT114), .ZN(n775) );
  NAND2_X1 U724 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  INV_X1 U725 ( .A(n691), .ZN(n654) );
  INV_X1 U726 ( .A(G952), .ZN(n656) );
  XNOR2_X1 U727 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT93), .B(KEYINPUT124), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT59), .ZN(n659) );
  XOR2_X1 U730 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n662) );
  NAND2_X1 U731 ( .A1(n397), .A2(G469), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n667), .A2(n749), .ZN(G54) );
  XNOR2_X1 U736 ( .A(n398), .B(n668), .ZN(G3) );
  NAND2_X1 U737 ( .A1(n683), .A2(n672), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT116), .ZN(n670) );
  XNOR2_X1 U739 ( .A(G104), .B(n670), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n674) );
  INV_X1 U741 ( .A(n671), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n672), .A2(n685), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G9) );
  XOR2_X1 U745 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n678) );
  NAND2_X1 U746 ( .A1(n681), .A2(n685), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U748 ( .A(G128), .B(n679), .ZN(G30) );
  XNOR2_X1 U749 ( .A(G143), .B(n680), .ZN(G45) );
  NAND2_X1 U750 ( .A1(n681), .A2(n683), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n682), .B(G146), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(G113), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(G116), .ZN(G18) );
  INV_X1 U756 ( .A(n764), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n690), .A2(KEYINPUT2), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n695) );
  INV_X1 U760 ( .A(n693), .ZN(n726) );
  NOR2_X1 U761 ( .A1(n726), .A2(n713), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n696), .A2(n765), .ZN(n734) );
  XNOR2_X1 U764 ( .A(KEYINPUT52), .B(KEYINPUT122), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n697), .B(KEYINPUT123), .ZN(n730) );
  NOR2_X1 U766 ( .A1(n539), .A2(n698), .ZN(n699) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n699), .Z(n700) );
  NOR2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U769 ( .A(KEYINPUT119), .B(n702), .Z(n708) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U771 ( .A(KEYINPUT50), .B(n705), .Z(n706) );
  XNOR2_X1 U772 ( .A(KEYINPUT120), .B(n706), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n711) );
  INV_X1 U774 ( .A(n709), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n712), .ZN(n714) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n728) );
  INV_X1 U778 ( .A(n715), .ZN(n717) );
  NAND2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n720), .B(KEYINPUT121), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U786 ( .A(n730), .B(n729), .Z(n731) );
  NOR2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U790 ( .A(n736), .Z(n739) );
  XOR2_X1 U791 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n737) );
  XNOR2_X1 U792 ( .A(n737), .B(KEYINPUT90), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n743), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U795 ( .A1(n397), .A2(G478), .ZN(n744) );
  NAND2_X1 U796 ( .A1(n397), .A2(G217), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U798 ( .A1(n749), .A2(n748), .ZN(G66) );
  NAND2_X1 U799 ( .A1(n750), .A2(n765), .ZN(n755) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U801 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n752), .A2(G898), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n753), .B(KEYINPUT126), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(n760) );
  XOR2_X1 U805 ( .A(n756), .B(n398), .Z(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U807 ( .A(n760), .B(n759), .Z(G69) );
  XNOR2_X1 U808 ( .A(n761), .B(KEYINPUT4), .ZN(n762) );
  XNOR2_X1 U809 ( .A(n763), .B(n762), .ZN(n767) );
  XNOR2_X1 U810 ( .A(n764), .B(n767), .ZN(n766) );
  NAND2_X1 U811 ( .A1(n766), .A2(n765), .ZN(n772) );
  XOR2_X1 U812 ( .A(G227), .B(n767), .Z(n768) );
  NAND2_X1 U813 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U814 ( .A1(G953), .A2(n769), .ZN(n770) );
  XOR2_X1 U815 ( .A(KEYINPUT127), .B(n770), .Z(n771) );
  NAND2_X1 U816 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U817 ( .A(G119), .B(n773), .Z(G21) );
  XOR2_X1 U818 ( .A(n774), .B(G131), .Z(G33) );
  XNOR2_X1 U819 ( .A(G134), .B(n775), .ZN(G36) );
  XOR2_X1 U820 ( .A(G137), .B(n776), .Z(G39) );
endmodule

