

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U547 ( .A(n517), .B(n516), .ZN(n874) );
  NOR2_X1 U548 ( .A1(G651), .A2(n624), .ZN(n650) );
  AND2_X1 U549 ( .A1(n512), .A2(G2104), .ZN(n875) );
  OR2_X1 U550 ( .A1(n764), .A2(n763), .ZN(n510) );
  AND2_X1 U551 ( .A1(n963), .A2(n809), .ZN(n511) );
  INV_X1 U552 ( .A(KEYINPUT26), .ZN(n687) );
  NOR2_X1 U553 ( .A1(n952), .A2(n691), .ZN(n697) );
  INV_X1 U554 ( .A(n726), .ZN(n711) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U556 ( .A(n710), .B(n709), .ZN(n715) );
  INV_X1 U557 ( .A(n956), .ZN(n745) );
  NOR2_X1 U558 ( .A1(n759), .A2(n745), .ZN(n746) );
  AND2_X1 U559 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U560 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n776) );
  NOR2_X1 U562 ( .A1(n797), .A2(n511), .ZN(n798) );
  XOR2_X1 U563 ( .A(KEYINPUT15), .B(n570), .Z(n820) );
  AND2_X1 U564 ( .A1(n521), .A2(n520), .ZN(G160) );
  INV_X1 U565 ( .A(G2105), .ZN(n512) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n512), .ZN(n879) );
  NAND2_X1 U567 ( .A1(n879), .A2(G125), .ZN(n515) );
  NAND2_X1 U568 ( .A1(G101), .A2(n875), .ZN(n513) );
  XOR2_X1 U569 ( .A(KEYINPUT23), .B(n513), .Z(n514) );
  AND2_X1 U570 ( .A1(n515), .A2(n514), .ZN(n521) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n517) );
  NOR2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NAND2_X1 U573 ( .A1(G137), .A2(n874), .ZN(n519) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U575 ( .A1(G113), .A2(n880), .ZN(n518) );
  AND2_X1 U576 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U577 ( .A1(G138), .A2(n874), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G102), .A2(n875), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n527) );
  NAND2_X1 U580 ( .A1(G126), .A2(n879), .ZN(n525) );
  NAND2_X1 U581 ( .A1(G114), .A2(n880), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n527), .A2(n526), .ZN(G164) );
  XNOR2_X1 U584 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U585 ( .A(KEYINPUT105), .B(G2435), .Z(n529) );
  XNOR2_X1 U586 ( .A(G2430), .B(G2438), .ZN(n528) );
  XNOR2_X1 U587 ( .A(n529), .B(n528), .ZN(n536) );
  XOR2_X1 U588 ( .A(G2446), .B(G2454), .Z(n531) );
  XNOR2_X1 U589 ( .A(G2451), .B(G2443), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U591 ( .A(n532), .B(G2427), .Z(n534) );
  XNOR2_X1 U592 ( .A(G1341), .B(G1348), .ZN(n533) );
  XNOR2_X1 U593 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U594 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U595 ( .A1(n537), .A2(G14), .ZN(G401) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n624) );
  INV_X1 U597 ( .A(G651), .ZN(n545) );
  NOR2_X1 U598 ( .A1(n624), .A2(n545), .ZN(n645) );
  NAND2_X1 U599 ( .A1(n645), .A2(G77), .ZN(n538) );
  XOR2_X1 U600 ( .A(KEYINPUT69), .B(n538), .Z(n541) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(KEYINPUT64), .ZN(n646) );
  NAND2_X1 U603 ( .A1(G90), .A2(n646), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(KEYINPUT9), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G52), .A2(n650), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n549) );
  NOR2_X1 U608 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X2 U609 ( .A(KEYINPUT1), .B(n546), .Z(n651) );
  NAND2_X1 U610 ( .A1(n651), .A2(G64), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT68), .B(n547), .Z(n548) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n814) );
  NAND2_X1 U617 ( .A1(n814), .A2(G567), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT11), .B(n551), .Z(G234) );
  NAND2_X1 U619 ( .A1(G56), .A2(n651), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n552), .Z(n559) );
  NAND2_X1 U621 ( .A1(n646), .A2(G81), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT75), .B(n553), .Z(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(KEYINPUT12), .ZN(n556) );
  NAND2_X1 U624 ( .A1(G68), .A2(n645), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n557), .Z(n558) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n650), .A2(G43), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n952) );
  INV_X1 U630 ( .A(G860), .ZN(n595) );
  OR2_X1 U631 ( .A1(n952), .A2(n595), .ZN(G153) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G79), .A2(n645), .ZN(n563) );
  NAND2_X1 U634 ( .A1(G54), .A2(n650), .ZN(n562) );
  NAND2_X1 U635 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n651), .A2(G66), .ZN(n564) );
  XNOR2_X1 U637 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U638 ( .A1(G92), .A2(n646), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U640 ( .A(KEYINPUT77), .B(n567), .Z(n568) );
  NOR2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U642 ( .A(n820), .ZN(n967) );
  NOR2_X1 U643 ( .A1(G868), .A2(n967), .ZN(n572) );
  INV_X1 U644 ( .A(G868), .ZN(n664) );
  NOR2_X1 U645 ( .A1(n664), .A2(G301), .ZN(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U647 ( .A(KEYINPUT78), .B(n573), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G51), .A2(n650), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G63), .A2(n651), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U651 ( .A(KEYINPUT6), .B(n576), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G89), .A2(n646), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n577), .B(KEYINPUT4), .ZN(n579) );
  NAND2_X1 U654 ( .A1(G76), .A2(n645), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U656 ( .A(n580), .B(KEYINPUT5), .Z(n581) );
  NOR2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U658 ( .A(KEYINPUT7), .B(n583), .Z(n585) );
  XOR2_X1 U659 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n584) );
  XNOR2_X1 U660 ( .A(n585), .B(n584), .ZN(G168) );
  XOR2_X1 U661 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U662 ( .A1(n645), .A2(G78), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G91), .A2(n646), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT70), .B(n588), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G53), .A2(n650), .ZN(n590) );
  NAND2_X1 U667 ( .A1(G65), .A2(n651), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n957) );
  XNOR2_X1 U670 ( .A(n957), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G299), .A2(n664), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n596), .A2(n820), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT16), .ZN(n598) );
  XOR2_X1 U677 ( .A(KEYINPUT81), .B(n598), .Z(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n952), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n820), .A2(G868), .ZN(n599) );
  NOR2_X1 U680 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n879), .ZN(n602) );
  XNOR2_X1 U683 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n875), .A2(G99), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G135), .A2(n874), .ZN(n606) );
  NAND2_X1 U687 ( .A1(G111), .A2(n880), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n899) );
  XOR2_X1 U690 ( .A(n899), .B(G2096), .Z(n609) );
  NOR2_X1 U691 ( .A1(G2100), .A2(n609), .ZN(n610) );
  XOR2_X1 U692 ( .A(KEYINPUT82), .B(n610), .Z(G156) );
  NAND2_X1 U693 ( .A1(n651), .A2(G67), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G93), .A2(n646), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G80), .A2(n645), .ZN(n614) );
  NAND2_X1 U697 ( .A1(G55), .A2(n650), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n665) );
  XNOR2_X1 U700 ( .A(n952), .B(KEYINPUT83), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n820), .A2(G559), .ZN(n617) );
  XNOR2_X1 U702 ( .A(n618), .B(n617), .ZN(n662) );
  XOR2_X1 U703 ( .A(n662), .B(KEYINPUT84), .Z(n619) );
  NOR2_X1 U704 ( .A1(G860), .A2(n619), .ZN(n620) );
  XOR2_X1 U705 ( .A(n665), .B(n620), .Z(G145) );
  NAND2_X1 U706 ( .A1(G49), .A2(n650), .ZN(n622) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U709 ( .A1(n651), .A2(n623), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G87), .A2(n624), .ZN(n625) );
  XOR2_X1 U711 ( .A(KEYINPUT85), .B(n625), .Z(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(n628), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G73), .A2(n645), .ZN(n629) );
  XNOR2_X1 U715 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n651), .A2(G61), .ZN(n631) );
  NAND2_X1 U717 ( .A1(G86), .A2(n646), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U719 ( .A1(G48), .A2(n650), .ZN(n632) );
  XNOR2_X1 U720 ( .A(KEYINPUT87), .B(n632), .ZN(n633) );
  NOR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G72), .A2(n645), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G47), .A2(n650), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n646), .A2(G85), .ZN(n639) );
  XOR2_X1 U727 ( .A(KEYINPUT66), .B(n639), .Z(n640) );
  NOR2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n651), .A2(G60), .ZN(n642) );
  XOR2_X1 U730 ( .A(KEYINPUT67), .B(n642), .Z(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(G290) );
  NAND2_X1 U732 ( .A1(n645), .A2(G75), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G88), .A2(n646), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U735 ( .A(KEYINPUT89), .B(n649), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G50), .A2(n650), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G62), .A2(n651), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U739 ( .A(KEYINPUT88), .B(n654), .Z(n655) );
  NAND2_X1 U740 ( .A1(n656), .A2(n655), .ZN(G303) );
  INV_X1 U741 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(n665), .ZN(n657) );
  XNOR2_X1 U743 ( .A(G305), .B(n657), .ZN(n658) );
  XNOR2_X1 U744 ( .A(G288), .B(n658), .ZN(n660) );
  XNOR2_X1 U745 ( .A(G290), .B(G166), .ZN(n659) );
  XNOR2_X1 U746 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n661), .B(G299), .ZN(n823) );
  XOR2_X1 U748 ( .A(n823), .B(n662), .Z(n663) );
  NOR2_X1 U749 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U750 ( .A1(G868), .A2(n665), .ZN(n666) );
  NOR2_X1 U751 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U754 ( .A1(n669), .A2(G2090), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n670), .B(KEYINPUT21), .ZN(n671) );
  XNOR2_X1 U756 ( .A(KEYINPUT90), .B(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n672), .ZN(G158) );
  XOR2_X1 U758 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XOR2_X1 U759 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U760 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U762 ( .A1(G237), .A2(n673), .ZN(n674) );
  XNOR2_X1 U763 ( .A(KEYINPUT92), .B(n674), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n675), .A2(G108), .ZN(n818) );
  NAND2_X1 U765 ( .A1(G567), .A2(n818), .ZN(n676) );
  XNOR2_X1 U766 ( .A(n676), .B(KEYINPUT93), .ZN(n682) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U768 ( .A(KEYINPUT91), .B(n677), .Z(n678) );
  XNOR2_X1 U769 ( .A(KEYINPUT22), .B(n678), .ZN(n679) );
  NAND2_X1 U770 ( .A1(n679), .A2(G96), .ZN(n680) );
  OR2_X1 U771 ( .A1(G218), .A2(n680), .ZN(n819) );
  AND2_X1 U772 ( .A1(G2106), .A2(n819), .ZN(n681) );
  NOR2_X1 U773 ( .A1(n682), .A2(n681), .ZN(G319) );
  INV_X1 U774 ( .A(G319), .ZN(n892) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U776 ( .A1(n892), .A2(n683), .ZN(n817) );
  NAND2_X1 U777 ( .A1(n817), .A2(G36), .ZN(G176) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n775) );
  INV_X1 U779 ( .A(n775), .ZN(n684) );
  NAND2_X1 U780 ( .A1(n776), .A2(n684), .ZN(n726) );
  NAND2_X1 U781 ( .A1(G8), .A2(n726), .ZN(n759) );
  NOR2_X1 U782 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XOR2_X1 U783 ( .A(n685), .B(KEYINPUT24), .Z(n686) );
  NOR2_X1 U784 ( .A1(n759), .A2(n686), .ZN(n764) );
  AND2_X1 U785 ( .A1(n711), .A2(G1996), .ZN(n688) );
  XNOR2_X1 U786 ( .A(n688), .B(n687), .ZN(n690) );
  NAND2_X1 U787 ( .A1(n726), .A2(G1341), .ZN(n689) );
  NAND2_X1 U788 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U789 ( .A1(n697), .A2(n820), .ZN(n695) );
  NOR2_X1 U790 ( .A1(n711), .A2(G1348), .ZN(n693) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n726), .ZN(n692) );
  NOR2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U793 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U794 ( .A(n696), .B(KEYINPUT98), .ZN(n699) );
  OR2_X1 U795 ( .A1(n697), .A2(n820), .ZN(n698) );
  NAND2_X1 U796 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n711), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U798 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U799 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U800 ( .A1(n975), .A2(n711), .ZN(n701) );
  NOR2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n957), .A2(n705), .ZN(n703) );
  NAND2_X1 U803 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n957), .A2(n705), .ZN(n706) );
  XOR2_X1 U805 ( .A(n706), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n710) );
  OR2_X1 U807 ( .A1(n711), .A2(G1961), .ZN(n713) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n932) );
  NAND2_X1 U809 ( .A1(n711), .A2(n932), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n716), .A2(G171), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n725) );
  NOR2_X1 U813 ( .A1(G171), .A2(n716), .ZN(n722) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n759), .ZN(n739) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n726), .ZN(n736) );
  NOR2_X1 U816 ( .A1(n739), .A2(n736), .ZN(n717) );
  NAND2_X1 U817 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n718), .ZN(n719) );
  XOR2_X1 U819 ( .A(KEYINPUT99), .B(n719), .Z(n720) );
  NOR2_X1 U820 ( .A1(n720), .A2(G168), .ZN(n721) );
  NOR2_X1 U821 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U823 ( .A1(n725), .A2(n724), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n737), .A2(G286), .ZN(n732) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n759), .ZN(n728) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U828 ( .A(n729), .B(KEYINPUT100), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n733), .A2(G8), .ZN(n735) );
  XOR2_X1 U832 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n734) );
  XNOR2_X1 U833 ( .A(n735), .B(n734), .ZN(n743) );
  NAND2_X1 U834 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U835 ( .A(n737), .ZN(n738) );
  NOR2_X1 U836 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U838 ( .A1(n743), .A2(n742), .ZN(n757) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U841 ( .A1(n749), .A2(n744), .ZN(n961) );
  NAND2_X1 U842 ( .A1(n757), .A2(n961), .ZN(n747) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n956) );
  NOR2_X1 U844 ( .A1(KEYINPUT33), .A2(n748), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U846 ( .A1(n750), .A2(n759), .ZN(n751) );
  XOR2_X1 U847 ( .A(G1981), .B(KEYINPUT102), .Z(n753) );
  XNOR2_X1 U848 ( .A(G305), .B(n753), .ZN(n949) );
  NAND2_X1 U849 ( .A1(n754), .A2(n949), .ZN(n762) );
  NAND2_X1 U850 ( .A1(G8), .A2(G166), .ZN(n755) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n755), .ZN(n756) );
  XNOR2_X1 U852 ( .A(n756), .B(KEYINPUT103), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U856 ( .A1(G140), .A2(n874), .ZN(n766) );
  NAND2_X1 U857 ( .A1(G104), .A2(n875), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n767), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n879), .A2(G128), .ZN(n768) );
  XNOR2_X1 U861 ( .A(n768), .B(KEYINPUT94), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G116), .A2(n880), .ZN(n769) );
  NAND2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n771), .Z(n772) );
  NOR2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U866 ( .A(KEYINPUT36), .B(n774), .ZN(n888) );
  XNOR2_X1 U867 ( .A(KEYINPUT37), .B(G2067), .ZN(n799) );
  NOR2_X1 U868 ( .A1(n888), .A2(n799), .ZN(n920) );
  NOR2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n809) );
  NAND2_X1 U870 ( .A1(n920), .A2(n809), .ZN(n777) );
  XOR2_X1 U871 ( .A(KEYINPUT95), .B(n777), .Z(n806) );
  NAND2_X1 U872 ( .A1(G131), .A2(n874), .ZN(n779) );
  NAND2_X1 U873 ( .A1(G95), .A2(n875), .ZN(n778) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G119), .A2(n879), .ZN(n781) );
  NAND2_X1 U876 ( .A1(G107), .A2(n880), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n855) );
  INV_X1 U879 ( .A(G1991), .ZN(n925) );
  NOR2_X1 U880 ( .A1(n855), .A2(n925), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G141), .A2(n874), .ZN(n784) );
  XNOR2_X1 U882 ( .A(n784), .B(KEYINPUT96), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G129), .A2(n879), .ZN(n786) );
  NAND2_X1 U884 ( .A1(G117), .A2(n880), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n875), .A2(G105), .ZN(n787) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U888 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n862) );
  AND2_X1 U890 ( .A1(n862), .A2(G1996), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n909) );
  INV_X1 U892 ( .A(n809), .ZN(n794) );
  NOR2_X1 U893 ( .A1(n909), .A2(n794), .ZN(n802) );
  INV_X1 U894 ( .A(n802), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n806), .A2(n795), .ZN(n796) );
  XOR2_X1 U896 ( .A(KEYINPUT97), .B(n796), .Z(n797) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n963) );
  NAND2_X1 U898 ( .A1(n510), .A2(n798), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n888), .A2(n799), .ZN(n917) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n862), .ZN(n904) );
  AND2_X1 U901 ( .A1(n925), .A2(n855), .ZN(n900) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U903 ( .A1(n900), .A2(n800), .ZN(n801) );
  NOR2_X1 U904 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U905 ( .A1(n904), .A2(n803), .ZN(n804) );
  XNOR2_X1 U906 ( .A(KEYINPUT104), .B(n804), .ZN(n805) );
  XNOR2_X1 U907 ( .A(n805), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U908 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U909 ( .A1(n917), .A2(n808), .ZN(n810) );
  NAND2_X1 U910 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U912 ( .A(KEYINPUT40), .B(n813), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n814), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n815) );
  NAND2_X1 U915 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U917 ( .A1(n817), .A2(n816), .ZN(G188) );
  NOR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(G325) );
  XOR2_X1 U919 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U925 ( .A(n952), .B(KEYINPUT116), .ZN(n822) );
  XNOR2_X1 U926 ( .A(G171), .B(n820), .ZN(n821) );
  XNOR2_X1 U927 ( .A(n822), .B(n821), .ZN(n825) );
  XOR2_X1 U928 ( .A(G286), .B(n823), .Z(n824) );
  XNOR2_X1 U929 ( .A(n825), .B(n824), .ZN(n826) );
  NOR2_X1 U930 ( .A1(G37), .A2(n826), .ZN(G397) );
  XNOR2_X1 U931 ( .A(G1966), .B(KEYINPUT41), .ZN(n836) );
  XOR2_X1 U932 ( .A(G1981), .B(G1971), .Z(n828) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1961), .ZN(n827) );
  XNOR2_X1 U934 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U935 ( .A(G1976), .B(G1956), .Z(n830) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U937 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U938 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U939 ( .A(KEYINPUT110), .B(G2474), .ZN(n833) );
  XNOR2_X1 U940 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n836), .B(n835), .ZN(G229) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2072), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n837), .B(G2678), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n839) );
  XNOR2_X1 U945 ( .A(KEYINPUT43), .B(G2096), .ZN(n838) );
  XNOR2_X1 U946 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U947 ( .A(G2100), .B(G2090), .Z(n841) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2084), .ZN(n840) );
  XNOR2_X1 U949 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U950 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U951 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n844) );
  XNOR2_X1 U952 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U953 ( .A(n847), .B(n846), .ZN(G227) );
  NAND2_X1 U954 ( .A1(G124), .A2(n879), .ZN(n848) );
  XNOR2_X1 U955 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U956 ( .A1(n875), .A2(G100), .ZN(n849) );
  NAND2_X1 U957 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G136), .A2(n874), .ZN(n852) );
  NAND2_X1 U959 ( .A1(G112), .A2(n880), .ZN(n851) );
  NAND2_X1 U960 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U961 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U962 ( .A(n899), .B(G162), .Z(n857) );
  XNOR2_X1 U963 ( .A(G160), .B(n855), .ZN(n856) );
  XNOR2_X1 U964 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n859) );
  XNOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n858) );
  XNOR2_X1 U967 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U968 ( .A(n861), .B(n860), .Z(n864) );
  XOR2_X1 U969 ( .A(G164), .B(n862), .Z(n863) );
  XNOR2_X1 U970 ( .A(n864), .B(n863), .ZN(n890) );
  NAND2_X1 U971 ( .A1(G118), .A2(n880), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n879), .A2(G130), .ZN(n865) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n865), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G142), .A2(n874), .ZN(n867) );
  NAND2_X1 U975 ( .A1(G106), .A2(n875), .ZN(n866) );
  NAND2_X1 U976 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U977 ( .A(KEYINPUT112), .B(n868), .Z(n869) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n869), .ZN(n870) );
  NOR2_X1 U979 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U980 ( .A1(n873), .A2(n872), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U982 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U983 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n878), .Z(n885) );
  NAND2_X1 U985 ( .A1(G127), .A2(n879), .ZN(n882) );
  NAND2_X1 U986 ( .A1(G115), .A2(n880), .ZN(n881) );
  NAND2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n910) );
  XNOR2_X1 U990 ( .A(n886), .B(n910), .ZN(n887) );
  XOR2_X1 U991 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U993 ( .A1(G37), .A2(n891), .ZN(G395) );
  NOR2_X1 U994 ( .A1(G401), .A2(n892), .ZN(n896) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n893) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n893), .ZN(n894) );
  NOR2_X1 U997 ( .A1(G397), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U999 ( .A1(n897), .A2(G395), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n898), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1002 ( .A(G160), .B(G2084), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n907) );
  XOR2_X1 U1005 ( .A(G2090), .B(G162), .Z(n903) );
  NOR2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n905), .B(KEYINPUT51), .ZN(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n916) );
  XOR2_X1 U1010 ( .A(G2072), .B(n910), .Z(n912) );
  XOR2_X1 U1011 ( .A(G164), .B(G2078), .Z(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1013 ( .A(KEYINPUT50), .B(n913), .Z(n914) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(n914), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT52), .B(n921), .ZN(n923) );
  INV_X1 U1019 ( .A(KEYINPUT55), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n924), .A2(G29), .ZN(n1004) );
  XNOR2_X1 U1022 ( .A(n925), .B(G25), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n926), .A2(G28), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT119), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G1996), .B(G32), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G2072), .B(G33), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G2067), .B(G26), .Z(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT120), .B(n932), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G27), .B(n933), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT53), .B(n938), .Z(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(G34), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G2084), .B(n940), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(n945), .Z(n946) );
  NOR2_X1 U1042 ( .A1(G29), .A2(n946), .ZN(n947) );
  XOR2_X1 U1043 ( .A(KEYINPUT122), .B(n947), .Z(n948) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n948), .ZN(n1002) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XNOR2_X1 U1046 ( .A(G168), .B(G1966), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(n951), .B(KEYINPUT57), .ZN(n971) );
  XNOR2_X1 U1049 ( .A(G301), .B(G1961), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n952), .B(G1341), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n966) );
  NAND2_X1 U1052 ( .A1(G1971), .A2(G303), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1054 ( .A(n957), .B(G1956), .Z(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT123), .B(n964), .Z(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(G1348), .B(n967), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n1000) );
  INV_X1 U1064 ( .A(G16), .ZN(n998) );
  XNOR2_X1 U1065 ( .A(KEYINPUT125), .B(G1966), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n974), .B(G21), .ZN(n993) );
  XNOR2_X1 U1067 ( .A(n975), .B(G20), .ZN(n983) );
  XOR2_X1 U1068 ( .A(G1341), .B(G19), .Z(n978) );
  XOR2_X1 U1069 ( .A(G6), .B(KEYINPUT124), .Z(n976) );
  XNOR2_X1 U1070 ( .A(G1981), .B(n976), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n979) );
  XNOR2_X1 U1073 ( .A(G4), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n984), .B(KEYINPUT60), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G5), .B(G1961), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT61), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1005), .B(KEYINPUT126), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT62), .B(n1006), .ZN(G150) );
  INV_X1 U1094 ( .A(G150), .ZN(G311) );
endmodule

