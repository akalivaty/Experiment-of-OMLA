//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1278, new_n1279, new_n1280, new_n1281;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  XNOR2_X1  g024(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G137), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(G2105), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n477), .A2(G136), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(KEYINPUT4), .A2(G138), .ZN(new_n484));
  OR2_X1    g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n462), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n485), .B2(new_n486), .ZN(new_n491));
  AND2_X1   g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G651), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G651), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(new_n502), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n511), .A2(G63), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n504), .A2(G89), .A3(new_n513), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n504), .A2(G51), .A3(G543), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G168));
  NAND3_X1  g100(.A1(new_n504), .A2(G52), .A3(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n504), .A2(G90), .A3(new_n513), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI211_X1 g105(.A(KEYINPUT72), .B(new_n529), .C1(new_n510), .C2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n510), .B2(new_n530), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n502), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n528), .B1(new_n531), .B2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n510), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n504), .A2(G81), .A3(new_n513), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n504), .A2(G43), .A3(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  XNOR2_X1  g125(.A(KEYINPUT77), .B(G65), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n513), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT76), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n504), .A2(G91), .A3(new_n513), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  AND2_X1   g134(.A1(G53), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n559), .B1(new_n504), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n504), .A2(new_n559), .A3(new_n560), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n556), .B(new_n557), .C1(new_n561), .C2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n534), .A2(new_n531), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n526), .A2(new_n527), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G301));
  NAND2_X1  g141(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n521), .A2(new_n568), .A3(new_n522), .A4(new_n523), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n567), .A2(new_n569), .ZN(G286));
  OR2_X1    g145(.A1(new_n507), .A2(new_n516), .ZN(G303));
  NAND3_X1  g146(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n504), .A2(G87), .A3(new_n513), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n513), .B2(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n576), .B1(new_n579), .B2(new_n502), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n501), .A2(new_n503), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n500), .A2(G651), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n581), .A2(G86), .A3(new_n582), .A4(new_n513), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n581), .A2(G48), .A3(G543), .A4(new_n582), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n508), .B2(new_n509), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(KEYINPUT79), .A3(G651), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n580), .A2(new_n583), .A3(new_n584), .A4(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT79), .B1(new_n586), .B2(G651), .ZN(new_n592));
  AOI211_X1 g167(.A(new_n576), .B(new_n502), .C1(new_n585), .C2(new_n577), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n583), .A2(new_n584), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n510), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n504), .A2(G85), .A3(new_n513), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n504), .A2(G47), .A3(G543), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G301), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n510), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n504), .A2(G54), .A3(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n514), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .A4(new_n513), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT81), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n608), .B1(new_n620), .B2(new_n607), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT82), .ZN(G284));
  XNOR2_X1  g197(.A(new_n621), .B(KEYINPUT83), .ZN(G321));
  AND2_X1   g198(.A1(G286), .A2(G868), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n556), .A2(new_n557), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n562), .A2(new_n561), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n629), .ZN(G297));
  OAI211_X1 g205(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n629), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n620), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n542), .A2(new_n607), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n620), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n477), .A2(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n477), .A2(G135), .ZN(new_n644));
  NOR2_X1   g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n473), .A2(G123), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT85), .B1(new_n473), .B2(G123), .ZN(new_n650));
  OAI221_X1 g225(.A(new_n644), .B1(new_n645), .B2(new_n646), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n642), .A2(new_n643), .A3(new_n653), .ZN(G156));
  INV_X1    g229(.A(G14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n657), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n663), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n656), .A3(new_n667), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT86), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n655), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n670), .A2(new_n672), .ZN(new_n678));
  AOI21_X1  g253(.A(KEYINPUT87), .B1(new_n678), .B2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n673), .A2(new_n680), .A3(new_n676), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G401));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT18), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(KEYINPUT18), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n686), .B(KEYINPUT89), .ZN(new_n693));
  INV_X1    g268(.A(new_n685), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n684), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n685), .B(KEYINPUT17), .Z(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n684), .A3(new_n693), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT90), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n690), .C2(new_n691), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n703), .A3(new_n652), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n652), .B1(new_n700), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n641), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(G2100), .A3(new_n704), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(G227));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  INV_X1    g286(.A(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1971), .B(G1976), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(G1956), .B(G2474), .Z(new_n718));
  XOR2_X1   g293(.A(G1961), .B(G1966), .Z(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT20), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n719), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n717), .A2(new_n720), .A3(new_n723), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G1986), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n721), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n724), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G1986), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n727), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(new_n727), .B2(new_n733), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n714), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n727), .A2(new_n733), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(new_n734), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n741), .A2(new_n713), .A3(new_n736), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(G229));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n477), .A2(G131), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n473), .A2(G119), .ZN(new_n747));
  OR2_X1    g322(.A1(G95), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n744), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  XOR2_X1   g328(.A(new_n752), .B(new_n753), .Z(new_n754));
  INV_X1    g329(.A(G290), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G16), .B2(G24), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(new_n732), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n732), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n754), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G16), .ZN(new_n763));
  NOR2_X1   g338(.A1(G166), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(G22), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n763), .A2(G23), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G288), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT33), .B(G1976), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n598), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G6), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n773), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n762), .B1(new_n779), .B2(KEYINPUT34), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT34), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n773), .A2(new_n777), .A3(new_n781), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(KEYINPUT36), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(KEYINPUT36), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n744), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n477), .A2(G140), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n473), .A2(G128), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT92), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n789), .B1(new_n800), .B2(new_n744), .ZN(new_n801));
  INV_X1    g376(.A(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n763), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n763), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n803), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n744), .A2(G32), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n477), .A2(G141), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n473), .A2(G129), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT26), .Z(new_n813));
  NAND3_X1  g388(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n810), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n809), .B1(new_n816), .B2(new_n744), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT27), .B(G1996), .Z(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  NAND2_X1  g394(.A1(G164), .A2(G29), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G27), .B2(G29), .ZN(new_n821));
  INV_X1    g396(.A(G2078), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n763), .A2(G21), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G168), .B2(new_n763), .ZN(new_n827));
  INV_X1    g402(.A(G1966), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n763), .A2(G19), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n543), .B2(new_n763), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G1341), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n832), .C1(G1961), .C2(new_n806), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n651), .A2(new_n744), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT30), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G28), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n744), .B1(new_n835), .B2(G28), .ZN(new_n837));
  AND2_X1   g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  NOR2_X1   g413(.A1(KEYINPUT31), .A2(G11), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n836), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n831), .A2(G1341), .ZN(new_n842));
  AND2_X1   g417(.A1(KEYINPUT24), .A2(G34), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n744), .B1(KEYINPUT24), .B2(G34), .ZN(new_n844));
  OAI22_X1  g419(.A1(G160), .A2(new_n744), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(G2084), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(G2084), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n841), .A2(new_n842), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NOR4_X1   g423(.A1(new_n808), .A2(new_n825), .A3(new_n833), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n744), .A2(G35), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G162), .B2(new_n744), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(new_n850), .C1(G162), .C2(new_n744), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n852), .A2(KEYINPUT29), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT29), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(G2090), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n763), .A2(G20), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n629), .B2(new_n763), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G1956), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT101), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n849), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT25), .ZN(new_n867));
  NAND2_X1  g442(.A1(G103), .A2(G2104), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(G2105), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n477), .A2(G139), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(G115), .A2(G2104), .ZN(new_n872));
  INV_X1    g447(.A(G127), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n472), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G2105), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT95), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(KEYINPUT96), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT96), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G29), .ZN(new_n883));
  NOR2_X1   g458(.A1(G29), .A2(G33), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT94), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G2072), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT98), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n763), .A2(G4), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n620), .B2(new_n763), .ZN(new_n891));
  INV_X1    g466(.A(G1348), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n886), .A2(KEYINPUT97), .A3(new_n887), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT97), .B1(new_n886), .B2(new_n887), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  INV_X1    g473(.A(new_n858), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n900));
  INV_X1    g475(.A(new_n863), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n866), .A2(new_n897), .A3(new_n898), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n902), .A2(new_n864), .A3(new_n865), .A4(new_n849), .ZN(new_n904));
  INV_X1    g479(.A(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT102), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n786), .A2(new_n787), .B1(new_n903), .B2(new_n906), .ZN(G311));
  AOI211_X1 g482(.A(new_n784), .B(KEYINPUT36), .C1(new_n780), .C2(new_n782), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n783), .A2(new_n785), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n787), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(G150));
  NAND3_X1  g487(.A1(new_n504), .A2(G93), .A3(new_n513), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n913), .B(new_n914), .C1(new_n502), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G860), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT37), .Z(new_n918));
  OR2_X1    g493(.A1(new_n916), .A2(new_n542), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n542), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n620), .A2(G559), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT103), .ZN(new_n927));
  INV_X1    g502(.A(G860), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n918), .B1(new_n927), .B2(new_n929), .ZN(G145));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n651), .B(G160), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G162), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n477), .A2(G142), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n473), .A2(G130), .ZN(new_n935));
  NOR2_X1   g510(.A1(G106), .A2(G2105), .ZN(new_n936));
  OAI21_X1  g511(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n639), .B(new_n938), .Z(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(new_n750), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n497), .A2(KEYINPUT104), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n489), .A2(new_n493), .A3(new_n942), .A4(new_n496), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n815), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n798), .A2(new_n799), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n792), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n815), .A3(new_n943), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n941), .A2(new_n815), .A3(new_n943), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n800), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n882), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n877), .A2(new_n879), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n933), .B1(new_n940), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n949), .A2(new_n951), .A3(new_n955), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n882), .B1(new_n949), .B2(new_n951), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n954), .A2(new_n962), .A3(new_n956), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n940), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI211_X1 g541(.A(KEYINPUT106), .B(new_n940), .C1(new_n961), .C2(new_n963), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n931), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n939), .B(new_n751), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT105), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n962), .B1(new_n954), .B2(new_n956), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n965), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(KEYINPUT107), .A3(new_n974), .A4(new_n958), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n969), .B1(new_n956), .B2(new_n954), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n957), .A2(new_n940), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n933), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT40), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT40), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n981), .C1(new_n968), .C2(new_n975), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(G395));
  OR2_X1    g561(.A1(new_n635), .A2(new_n921), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n617), .A2(new_n618), .ZN(new_n988));
  INV_X1    g563(.A(new_n614), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n629), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n619), .A2(G299), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n635), .A2(new_n921), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n987), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT41), .ZN(new_n996));
  INV_X1    g571(.A(new_n992), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n619), .A2(G299), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT41), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n987), .A2(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OR3_X1    g576(.A1(new_n995), .A2(new_n1001), .A3(KEYINPUT42), .ZN(new_n1002));
  OR2_X1    g577(.A1(G290), .A2(G288), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G290), .A2(G288), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT108), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n1006));
  AND2_X1   g581(.A1(G290), .A2(G288), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G290), .A2(G288), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G303), .B1(new_n590), .B2(new_n596), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G303), .A2(new_n590), .A3(new_n596), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1013), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1015), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT42), .B1(new_n995), .B2(new_n1001), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1002), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1002), .B2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g595(.A(G868), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n916), .A2(new_n607), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(G295));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1022), .ZN(G331));
  OR3_X1    g599(.A1(new_n1015), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1015), .A2(new_n1011), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n1010), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n999), .A2(new_n1000), .ZN(new_n1028));
  NAND3_X1  g603(.A1(G171), .A2(new_n567), .A3(new_n569), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G171), .A2(KEYINPUT109), .A3(new_n524), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(G301), .B2(G168), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n920), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n916), .A2(new_n542), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n919), .A2(new_n1037), .A3(new_n920), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT109), .B1(G171), .B2(new_n524), .ZN(new_n1041));
  NAND3_X1  g616(.A1(G301), .A2(G168), .A3(new_n1031), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(new_n1036), .A3(new_n1038), .A4(new_n1029), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1028), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1040), .A2(new_n1044), .B1(new_n992), .B2(new_n991), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1027), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1043), .A2(new_n1029), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n993), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1028), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1017), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n980), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT43), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT43), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1047), .A2(new_n1055), .A3(new_n1052), .A4(new_n980), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(KEYINPUT44), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1060));
  AOI21_X1  g635(.A(G37), .B1(new_n1060), .B2(new_n1027), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(KEYINPUT112), .A3(new_n1055), .A4(new_n1052), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1054), .A2(KEYINPUT111), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1053), .A2(new_n1065), .A3(KEYINPUT43), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(new_n1067), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g643(.A(G1384), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n941), .A2(new_n1069), .A3(new_n943), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT45), .ZN(new_n1071));
  AND2_X1   g646(.A1(G160), .A2(G40), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n800), .B(G2067), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n815), .B(G1996), .Z(new_n1076));
  OR2_X1    g651(.A1(new_n751), .A2(new_n753), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n751), .A2(new_n753), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G290), .B(G1986), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n497), .A2(new_n1069), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT50), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n497), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1082), .A2(new_n1084), .A3(new_n1072), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G160), .A2(G40), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1083), .B2(KEYINPUT50), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1082), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n892), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n497), .A2(G160), .A3(G40), .A4(new_n1069), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2067), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n990), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n628), .B2(KEYINPUT119), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n629), .ZN(new_n1098));
  OAI211_X1 g673(.A(G299), .B(new_n1096), .C1(KEYINPUT119), .C2(new_n628), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1084), .A2(new_n1072), .A3(new_n1086), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT118), .B(G1956), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1083), .A2(new_n1071), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT113), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1071), .A2(G1384), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n941), .A2(new_n943), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1069), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1105), .A2(new_n1072), .A3(new_n1107), .A4(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT56), .B(G2072), .Z(new_n1112));
  OAI211_X1 g687(.A(new_n1100), .B(new_n1103), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1095), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1112), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1072), .A3(new_n1105), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1100), .B1(new_n1118), .B2(new_n1103), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1101), .A2(KEYINPUT120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1089), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1348), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1123), .A2(new_n619), .A3(new_n1093), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1095), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1088), .A2(G1996), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1105), .A2(new_n1107), .A3(new_n1110), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1092), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1127), .A2(KEYINPUT121), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT121), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n543), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1113), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1119), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n543), .B(new_n1133), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1125), .A2(new_n1135), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1119), .A2(new_n1137), .A3(new_n1136), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1123), .A2(new_n1093), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1120), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1111), .B2(G2078), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n804), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n497), .A2(new_n1106), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1072), .A2(new_n1149), .ZN(new_n1150));
  OR4_X1    g725(.A1(new_n1146), .A2(new_n1150), .A3(G2078), .A4(new_n1108), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1088), .A2(new_n1146), .A3(G2078), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1107), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1147), .A2(new_n1148), .A3(G301), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n828), .B1(new_n1150), .B2(new_n1108), .ZN(new_n1161));
  INV_X1    g736(.A(G2084), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1084), .A2(new_n1162), .A3(new_n1072), .A4(new_n1086), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1160), .B(G8), .C1(new_n1164), .C2(new_n524), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n524), .A2(G8), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g744(.A(KEYINPUT123), .B(new_n1167), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1165), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1164), .A2(G8), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(KEYINPUT51), .A3(new_n1167), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1158), .A2(new_n1159), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT114), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(G303), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT55), .ZN(new_n1180));
  INV_X1    g755(.A(G8), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(G166), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1101), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1111), .A2(new_n766), .B1(new_n1185), .B2(new_n857), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1186), .B2(new_n1181), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1111), .A2(new_n766), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1101), .A2(G2090), .ZN(new_n1189));
  OAI211_X1 g764(.A(G8), .B(new_n1183), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n572), .A2(new_n573), .A3(G1976), .A4(new_n574), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1092), .A2(G8), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT52), .ZN(new_n1193));
  INV_X1    g768(.A(G1976), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT52), .B1(G288), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1195), .A2(new_n1092), .A3(G8), .A4(new_n1191), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1092), .A2(G8), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n588), .A2(G1981), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT115), .B(G1981), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n595), .A2(new_n580), .A3(new_n587), .A4(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1199), .A2(KEYINPUT49), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT49), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT116), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1198), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT49), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1202), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n712), .B1(new_n594), .B2(new_n595), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1210), .A2(KEYINPUT116), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1197), .B(KEYINPUT117), .C1(new_n1206), .C2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(KEYINPUT116), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1203), .A2(new_n1198), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT117), .B1(new_n1217), .B2(new_n1197), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1187), .B(new_n1190), .C1(new_n1213), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1197), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT117), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1212), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1225), .A2(KEYINPUT124), .A3(new_n1187), .A4(new_n1190), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1147), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1159), .B1(new_n1227), .B2(G171), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(G171), .B2(new_n1152), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1175), .A2(new_n1221), .A3(new_n1226), .A4(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1145), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g806(.A(new_n1174), .B(new_n1165), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1232));
  OR2_X1    g807(.A1(new_n1232), .A2(KEYINPUT62), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1153), .B1(new_n1232), .B2(KEYINPUT62), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1221), .A2(new_n1233), .A3(new_n1226), .A4(new_n1234), .ZN(new_n1235));
  OR3_X1    g810(.A1(new_n1222), .A2(G286), .A3(new_n1173), .ZN(new_n1236));
  INV_X1    g811(.A(new_n1187), .ZN(new_n1237));
  OAI21_X1  g812(.A(KEYINPUT63), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(new_n1222), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1190), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1217), .ZN(new_n1241));
  OR2_X1    g816(.A1(G288), .A2(G1976), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1202), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI22_X1  g818(.A1(new_n1239), .A2(new_n1240), .B1(new_n1243), .B2(new_n1198), .ZN(new_n1244));
  AND2_X1   g819(.A1(new_n1238), .A2(new_n1244), .ZN(new_n1245));
  NOR3_X1   g820(.A1(new_n1173), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1246));
  NAND4_X1  g821(.A1(new_n1225), .A2(new_n1246), .A3(new_n1187), .A4(new_n1190), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1235), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1081), .B1(new_n1231), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1079), .A2(new_n1074), .ZN(new_n1250));
  NAND3_X1  g825(.A1(new_n1074), .A2(new_n732), .A3(new_n755), .ZN(new_n1251));
  XNOR2_X1  g826(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OR2_X1    g828(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1254));
  NAND3_X1  g829(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1256));
  OAI22_X1  g831(.A1(new_n1256), .A2(new_n1078), .B1(G2067), .B2(new_n947), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1257), .A2(new_n1074), .ZN(new_n1258));
  INV_X1    g833(.A(KEYINPUT46), .ZN(new_n1259));
  OAI211_X1 g834(.A(new_n1075), .B(new_n816), .C1(new_n1259), .C2(G1996), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1259), .B1(new_n1073), .B2(G1996), .ZN(new_n1261));
  AOI22_X1  g836(.A1(new_n1260), .A2(new_n1074), .B1(KEYINPUT125), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g837(.A(new_n1262), .B1(KEYINPUT125), .B2(new_n1261), .ZN(new_n1263));
  INV_X1    g838(.A(KEYINPUT47), .ZN(new_n1264));
  OAI211_X1 g839(.A(new_n1255), .B(new_n1258), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g840(.A(new_n1265), .B1(new_n1264), .B2(new_n1263), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1249), .A2(new_n1266), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g842(.A(new_n981), .B1(new_n968), .B2(new_n975), .ZN(new_n1269));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1270));
  AOI21_X1  g844(.A(new_n460), .B1(new_n739), .B2(new_n742), .ZN(new_n1271));
  NAND2_X1  g845(.A1(new_n1271), .A2(new_n682), .ZN(new_n1272));
  OAI21_X1  g846(.A(new_n1270), .B1(new_n1272), .B2(G227), .ZN(new_n1273));
  INV_X1    g847(.A(G227), .ZN(new_n1274));
  NAND4_X1  g848(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n682), .A4(new_n1271), .ZN(new_n1275));
  AND2_X1   g849(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  NOR3_X1   g850(.A1(new_n1067), .A2(new_n1269), .A3(new_n1276), .ZN(G308));
  NAND2_X1  g851(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1278));
  NAND3_X1  g852(.A1(new_n1278), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1279));
  INV_X1    g853(.A(new_n1269), .ZN(new_n1280));
  NAND2_X1  g854(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1281));
  NAND3_X1  g855(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(G225));
endmodule


