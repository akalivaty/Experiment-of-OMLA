//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n208), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n232), .B(new_n235), .C1(new_n222), .C2(new_n223), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n225), .A2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n210), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT66), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G223), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n259), .B1(new_n216), .B2(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n264), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n229), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  INV_X1    g0080(.A(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT68), .B(G58), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n230), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n278), .B1(new_n267), .B2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(G50), .B2(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n276), .A2(G169), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(KEYINPUT69), .B1(new_n297), .B2(new_n276), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(KEYINPUT69), .B2(new_n296), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT70), .Z(new_n300));
  OR2_X1    g0100(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n211), .B1(new_n272), .B2(KEYINPUT71), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n271), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n265), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n308), .A3(KEYINPUT13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G169), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n311), .A2(new_n315), .A3(G169), .A4(new_n312), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n303), .A2(new_n308), .B1(new_n318), .B2(KEYINPUT13), .ZN(new_n319));
  OAI21_X1  g0119(.A(G179), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n210), .A2(G20), .ZN(new_n322));
  INV_X1    g0122(.A(new_n289), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n322), .B1(new_n286), .B2(new_n216), .C1(new_n323), .C2(new_n202), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n278), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT11), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(KEYINPUT73), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n267), .A2(G13), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n333), .B(new_n322), .C1(KEYINPUT74), .C2(KEYINPUT12), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n292), .A2(G68), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n331), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n321), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n291), .A2(new_n295), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(KEYINPUT9), .B1(new_n275), .B2(G200), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n276), .A2(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(KEYINPUT9), .C2(new_n342), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n292), .A2(G77), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G77), .B2(new_n294), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT8), .B(G58), .Z(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n287), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n279), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(new_n218), .B2(new_n257), .C1(new_n260), .C2(new_n211), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n265), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n271), .B1(G244), .B2(new_n273), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n362), .B2(G190), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n356), .B1(new_n362), .B2(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n361), .A2(G179), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n346), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G190), .B1(new_n317), .B2(new_n319), .ZN(new_n370));
  INV_X1    g0170(.A(new_n340), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n311), .A2(G200), .A3(new_n312), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n300), .A2(new_n341), .A3(new_n369), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  OR2_X1    g0177(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g0179(.A(G33), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G33), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n377), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n257), .B2(G20), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n210), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT68), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G58), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n201), .B1(new_n394), .B2(G68), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n395), .A2(new_n230), .B1(new_n396), .B2(new_n323), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n375), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n378), .A2(new_n400), .A3(G33), .A4(new_n379), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g0203(.A(G33), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(KEYINPUT3), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT76), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n230), .B(new_n401), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n378), .A2(G33), .A3(new_n379), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n400), .B1(KEYINPUT3), .B2(new_n404), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(new_n230), .A3(new_n388), .A4(new_n401), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(G68), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n397), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT79), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n375), .C1(new_n390), .C2(new_n397), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n399), .A2(new_n416), .A3(new_n278), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n284), .A2(new_n294), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n284), .B2(new_n292), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G169), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n401), .B1(new_n405), .B2(new_n407), .ZN(new_n424));
  NOR2_X1   g0224(.A1(G223), .A2(G1698), .ZN(new_n425));
  INV_X1    g0225(.A(G226), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n404), .A2(new_n212), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n264), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n264), .A2(G232), .A3(new_n268), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n270), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n423), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n427), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n412), .B2(new_n401), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n265), .B1(new_n436), .B2(new_n429), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n270), .A2(new_n432), .A3(KEYINPUT80), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT80), .B1(new_n270), .B2(new_n432), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n440), .A3(new_n297), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n422), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n442), .B1(new_n419), .B2(new_n421), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n364), .B1(new_n431), .B2(new_n433), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(new_n440), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n419), .A2(new_n421), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n419), .A2(KEYINPUT17), .A3(new_n452), .A4(new_n421), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n445), .A2(new_n448), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n374), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n424), .A2(KEYINPUT22), .A3(new_n230), .A4(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n212), .A2(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT22), .B1(new_n257), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n218), .A2(KEYINPUT23), .A3(G20), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT23), .B1(new_n218), .B2(G20), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n463), .A2(new_n464), .B1(G20), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n459), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n459), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n278), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n279), .B(new_n294), .C1(G1), .C2(new_n404), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n218), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n294), .ZN(new_n475));
  INV_X1    g0275(.A(new_n294), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n476), .A2(KEYINPUT87), .A3(KEYINPUT25), .A4(new_n218), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n472), .A2(G107), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G41), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n267), .B(G45), .C1(new_n480), .C2(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g0282(.A(G274), .ZN(new_n483));
  INV_X1    g0283(.A(new_n229), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n263), .ZN(new_n485));
  INV_X1    g0285(.A(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G41), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n482), .A2(new_n485), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n481), .B2(KEYINPUT82), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n495));
  OAI211_X1 g0295(.A(G264), .B(new_n264), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G294), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n404), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G250), .A2(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(G257), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G1698), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n424), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n493), .B(new_n496), .C1(new_n502), .C2(new_n264), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(KEYINPUT88), .A3(G169), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n297), .B2(new_n503), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT88), .B1(new_n503), .B2(G169), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n479), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n503), .A2(new_n364), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n503), .A2(G190), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n470), .B(new_n478), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n476), .A2(KEYINPUT84), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n294), .B2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n471), .B2(new_n512), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(G33), .B2(G283), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT81), .B(G97), .Z(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G33), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(G20), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT85), .B1(new_n278), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n278), .A2(KEYINPUT85), .A3(new_n521), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n520), .B(KEYINPUT20), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G257), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n219), .B2(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n424), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(G303), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n257), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n264), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G270), .B(new_n264), .C1(new_n494), .C2(new_n495), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n493), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT21), .B(G169), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n537), .ZN(new_n539));
  INV_X1    g0339(.A(new_n530), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n412), .B2(new_n401), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n265), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n542), .A3(G179), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n528), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n535), .B2(new_n537), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n539), .A2(new_n542), .A3(G190), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n528), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  OAI21_X1  g0349(.A(G169), .B1(new_n535), .B2(new_n537), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n528), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT86), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT86), .B(new_n549), .C1(new_n550), .C2(new_n528), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n544), .B(new_n548), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n424), .A2(new_n230), .A3(G68), .ZN(new_n556));
  OR2_X1    g0356(.A1(KEYINPUT81), .A2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT81), .A2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT19), .B1(new_n559), .B2(new_n287), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n519), .A2(new_n212), .A3(new_n218), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n230), .B1(new_n306), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n278), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n472), .A2(new_n352), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n351), .A2(new_n476), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G238), .A2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n217), .B2(G1698), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n412), .B2(new_n401), .ZN(new_n573));
  INV_X1    g0373(.A(new_n465), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n265), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n264), .B(G250), .C1(G1), .C2(new_n486), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n485), .A2(KEYINPUT83), .A3(new_n487), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n264), .A2(G274), .A3(new_n487), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n577), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n423), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n297), .A3(new_n582), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n569), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n264), .C1(new_n494), .C2(new_n495), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n493), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n217), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(new_n258), .A3(new_n406), .A4(new_n382), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n406), .A2(new_n382), .A3(G250), .A4(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n258), .A2(G244), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n424), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n589), .B(new_n297), .C1(new_n599), .C2(new_n264), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n218), .B1(new_n384), .B2(new_n389), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT6), .B1(new_n206), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n218), .A2(KEYINPUT6), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n557), .B2(new_n558), .ZN(new_n605));
  OAI21_X1  g0405(.A(G20), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n289), .A2(G77), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n278), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G97), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n476), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n471), .B2(new_n610), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n595), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n596), .B1(new_n412), .B2(new_n401), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(KEYINPUT4), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n588), .B1(new_n617), .B2(new_n265), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n600), .B(new_n614), .C1(G169), .C2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n589), .B(G190), .C1(new_n599), .C2(new_n264), .ZN(new_n620));
  INV_X1    g0420(.A(new_n377), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n404), .B1(new_n402), .B2(new_n403), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n382), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n385), .A2(new_n387), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n406), .A2(new_n382), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n230), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G107), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n607), .A3(new_n606), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n612), .B1(new_n628), .B2(new_n278), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n620), .B(new_n629), .C1(new_n364), .C2(new_n618), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n583), .A2(G200), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n565), .A2(new_n278), .B1(new_n476), .B2(new_n351), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n472), .A2(G87), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n575), .A2(G190), .A3(new_n582), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n586), .A2(new_n619), .A3(new_n630), .A4(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n458), .A2(new_n511), .A3(new_n555), .A4(new_n636), .ZN(G372));
  AND3_X1   g0437(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n341), .B1(new_n638), .B2(new_n368), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n455), .A2(new_n456), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n446), .A2(new_n447), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT18), .B(new_n442), .C1(new_n419), .C2(new_n421), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n346), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n458), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n583), .B2(new_n423), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT89), .B(G169), .C1(new_n575), .C2(new_n582), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n585), .B(new_n569), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n553), .A2(new_n554), .ZN(new_n653));
  INV_X1    g0453(.A(new_n544), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n507), .A3(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n510), .A2(new_n635), .A3(new_n619), .A4(new_n630), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n586), .A2(new_n635), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n658), .B2(new_n619), .ZN(new_n659));
  INV_X1    g0459(.A(new_n619), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n651), .A3(new_n661), .A4(new_n635), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n300), .B(new_n646), .C1(new_n647), .C2(new_n664), .ZN(G369));
  NAND2_X1  g0465(.A1(new_n653), .A2(new_n654), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n333), .A2(KEYINPUT27), .A3(G20), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT27), .B1(new_n333), .B2(G20), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n528), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n544), .B1(new_n553), .B2(new_n554), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n547), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n674), .B(new_n675), .C1(new_n677), .C2(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n479), .A2(new_n671), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n511), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n507), .A2(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n666), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n678), .A2(new_n682), .A3(G330), .A4(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n507), .A2(new_n671), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n507), .A2(new_n510), .A3(new_n672), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n666), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n561), .A2(G116), .ZN(new_n689));
  INV_X1    g0489(.A(new_n233), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n227), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n619), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n660), .A2(new_n651), .A3(new_n635), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(KEYINPUT26), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n671), .B1(new_n698), .B2(new_n657), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT93), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n671), .B1(new_n657), .B2(new_n663), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n700), .B(KEYINPUT93), .C1(KEYINPUT29), .C2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n686), .A2(new_n555), .A3(new_n636), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n671), .A2(KEYINPUT31), .ZN(new_n705));
  INV_X1    g0505(.A(new_n496), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n424), .A2(new_n501), .ZN(new_n707));
  INV_X1    g0507(.A(new_n498), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n265), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n579), .A2(new_n580), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT83), .B1(new_n485), .B2(new_n487), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n576), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n424), .A2(new_n571), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n465), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(new_n715), .B2(new_n265), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n618), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT91), .B1(new_n717), .B2(new_n543), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(new_n543), .ZN(new_n720));
  INV_X1    g0520(.A(new_n501), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n412), .B2(new_n401), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n265), .B1(new_n722), .B2(new_n498), .ZN(new_n723));
  AND4_X1   g0523(.A1(new_n723), .A2(new_n575), .A3(new_n496), .A4(new_n582), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n720), .A2(new_n724), .A3(new_n725), .A4(new_n618), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n718), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n720), .A2(new_n724), .A3(KEYINPUT30), .A4(new_n618), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n589), .B1(new_n599), .B2(new_n264), .ZN(new_n729));
  AOI21_X1  g0529(.A(G179), .B1(new_n575), .B2(new_n582), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n539), .A2(new_n542), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n503), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n705), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n730), .A2(new_n731), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT92), .A3(new_n503), .A4(new_n729), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT92), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n736), .A2(new_n738), .A3(new_n728), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n718), .A2(new_n719), .A3(new_n726), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n672), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n704), .B(new_n734), .C1(new_n741), .C2(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n701), .A2(new_n703), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n695), .B1(new_n744), .B2(G1), .ZN(G364));
  NAND3_X1  g0545(.A1(new_n678), .A2(G330), .A3(new_n683), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n230), .A2(G13), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n267), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n691), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n678), .A2(new_n683), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n230), .B1(KEYINPUT96), .B2(new_n423), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n423), .A2(KEYINPUT96), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n229), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n230), .A2(new_n297), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n450), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n230), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n450), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G50), .B1(new_n769), .B2(G107), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n450), .A2(G179), .A3(G200), .ZN(new_n771));
  OAI21_X1  g0571(.A(G97), .B1(new_n771), .B2(new_n230), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n765), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n770), .B(new_n772), .C1(new_n210), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(KEYINPUT32), .A3(new_n396), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT32), .B1(new_n777), .B2(new_n396), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n212), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n764), .A2(new_n776), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n764), .A2(G190), .A3(new_n364), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n257), .B1(new_n782), .B2(new_n216), .C1(new_n283), .C2(new_n783), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n775), .A2(new_n778), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n773), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G326), .ZN(new_n790));
  INV_X1    g0590(.A(new_n766), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n532), .B2(new_n780), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n783), .ZN(new_n793));
  INV_X1    g0593(.A(new_n777), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(G322), .B1(new_n794), .B2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n625), .C1(new_n796), .C2(new_n782), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n771), .A2(new_n230), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(new_n497), .B1(new_n768), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n792), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n763), .B1(new_n785), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n758), .A2(new_n763), .ZN(new_n803));
  INV_X1    g0603(.A(new_n424), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n233), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n250), .A2(new_n486), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n486), .C2(new_n228), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n257), .A2(new_n233), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(G116), .B2(new_n233), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n803), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n802), .A2(new_n812), .A3(new_n750), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n752), .A2(new_n755), .B1(new_n760), .B2(new_n813), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n368), .A2(new_n671), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n365), .B1(new_n355), .B2(new_n672), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n368), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n702), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n750), .B1(new_n818), .B2(new_n743), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n743), .B2(new_n818), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n799), .A2(new_n774), .B1(new_n791), .B2(new_n532), .ZN(new_n821));
  INV_X1    g0621(.A(new_n780), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G107), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n783), .A2(new_n497), .B1(new_n777), .B2(new_n796), .ZN(new_n824));
  INV_X1    g0624(.A(new_n782), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n257), .B(new_n824), .C1(G116), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n769), .A2(G87), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n772), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n793), .A2(G143), .B1(new_n825), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n791), .B2(new_n830), .C1(new_n831), .C2(new_n774), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n798), .A2(new_n283), .B1(new_n768), .B2(new_n210), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n780), .A2(new_n202), .B1(new_n777), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n804), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n832), .A2(new_n833), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n828), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n763), .ZN(new_n842));
  INV_X1    g0642(.A(new_n757), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n763), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n751), .B1(new_n844), .B2(new_n216), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n842), .B(new_n845), .C1(new_n817), .C2(new_n757), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n820), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  OR2_X1    g0648(.A1(new_n603), .A2(new_n605), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n851), .A4(new_n231), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI211_X1 g0653(.A(new_n228), .B(G77), .C1(new_n210), .C2(new_n283), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n267), .B(G13), .C1(new_n854), .C2(new_n246), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n421), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n210), .B1(new_n408), .B2(KEYINPUT7), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n397), .B1(new_n858), .B2(new_n413), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n279), .B1(new_n859), .B2(KEYINPUT16), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n414), .A2(new_n415), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n375), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n857), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT98), .B1(new_n863), .B2(new_n669), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n416), .A2(new_n278), .ZN(new_n865));
  INV_X1    g0665(.A(new_n375), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n421), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT98), .ZN(new_n869));
  INV_X1    g0669(.A(new_n669), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n443), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n453), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n419), .A2(new_n421), .A3(new_n452), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n446), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n422), .A2(new_n870), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n457), .A2(new_n872), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n815), .B1(new_n702), .B2(new_n817), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n340), .A2(new_n671), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n341), .A2(new_n373), .A3(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n340), .B(new_n671), .C1(new_n638), .C2(new_n321), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT97), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT97), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n341), .A2(new_n894), .A3(new_n373), .A4(new_n890), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n645), .A2(new_n669), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT99), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n902));
  AND4_X1   g0702(.A1(new_n878), .A2(new_n444), .A3(new_n879), .A4(new_n453), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n879), .B1(new_n644), .B2(new_n640), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n884), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n886), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT101), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n881), .B2(new_n882), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT101), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n906), .A2(new_n886), .A3(new_n913), .A4(new_n907), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n341), .A2(new_n671), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n897), .A2(KEYINPUT99), .A3(new_n898), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n901), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n646), .A2(new_n300), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n701), .A2(new_n703), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n458), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n919), .B(new_n922), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n886), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n736), .A2(new_n738), .A3(new_n728), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n705), .B1(new_n727), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n636), .A2(new_n676), .A3(new_n547), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n507), .A2(new_n510), .A3(new_n672), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n740), .A2(new_n738), .A3(new_n736), .A4(new_n728), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT31), .B1(new_n930), .B2(new_n671), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n893), .A2(new_n817), .A3(new_n895), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT40), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n935), .A2(KEYINPUT40), .B1(new_n887), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n647), .B2(new_n932), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n704), .B(new_n926), .C1(new_n741), .C2(KEYINPUT31), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n887), .A2(new_n936), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n924), .B2(new_n934), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n458), .B(new_n939), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n943), .A3(G330), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n923), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n267), .B2(new_n747), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n923), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n856), .B1(new_n946), .B2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n651), .A2(new_n635), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT102), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n672), .B1(new_n632), .B2(new_n633), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n652), .A2(new_n951), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n759), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n805), .A2(new_n244), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n803), .B1(new_n233), .B2(new_n351), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n750), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n774), .A2(new_n396), .B1(new_n210), .B2(new_n798), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n769), .A2(G77), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n791), .B2(new_n962), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n257), .B1(new_n782), .B2(new_n202), .C1(new_n831), .C2(new_n783), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n780), .A2(new_n283), .B1(new_n777), .B2(new_n830), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT106), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n780), .A2(new_n512), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT46), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n825), .A2(G283), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n793), .A2(G303), .B1(new_n794), .B2(G317), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n969), .A2(new_n804), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n766), .A2(G311), .B1(new_n769), .B2(new_n559), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n218), .B2(new_n798), .C1(new_n497), .C2(new_n774), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n965), .A2(new_n967), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n959), .B1(new_n976), .B2(new_n763), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n956), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n684), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n660), .A2(new_n671), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n619), .B(new_n630), .C1(new_n629), .C2(new_n672), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n687), .A2(new_n685), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n687), .A2(new_n982), .A3(KEYINPUT45), .A4(new_n685), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n982), .B1(new_n687), .B2(new_n685), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT44), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n991), .B(new_n982), .C1(new_n687), .C2(new_n685), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n979), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n987), .B(new_n684), .C1(new_n990), .C2(new_n992), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n676), .A2(new_n671), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n687), .B1(new_n682), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT105), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n746), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n746), .A2(new_n999), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n998), .B2(new_n1000), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n744), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n691), .B(KEYINPUT41), .Z(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n749), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n982), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n684), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT42), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n687), .B2(new_n1008), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n686), .A2(KEYINPUT42), .A3(new_n666), .A4(new_n982), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n619), .B1(new_n981), .B2(new_n507), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT103), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT103), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n619), .C1(new_n981), .C2(new_n507), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n672), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1013), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT104), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n955), .B(KEYINPUT43), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1009), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1009), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n978), .B1(new_n1007), .B2(new_n1028), .ZN(G387));
  NAND3_X1  g0829(.A1(new_n701), .A2(new_n703), .A3(new_n743), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1003), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n998), .B1(new_n746), .B2(new_n999), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n746), .B(new_n999), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(new_n1033), .B2(new_n998), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n744), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1035), .A3(new_n691), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n680), .A2(new_n681), .A3(new_n758), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n809), .A2(new_n689), .B1(G107), .B2(new_n233), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n241), .A2(new_n486), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT107), .Z(new_n1040));
  INV_X1    g0840(.A(new_n689), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n1041), .C1(G68), .C2(G77), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n349), .A2(new_n202), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT50), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n805), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1038), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n803), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n750), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n798), .A2(new_n351), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n791), .A2(new_n396), .B1(new_n780), .B2(new_n216), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G97), .C2(new_n769), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n285), .A2(new_n773), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT108), .B(G150), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n783), .A2(new_n202), .B1(new_n1053), .B2(new_n777), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n825), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n424), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n798), .A2(new_n799), .B1(new_n780), .B2(new_n497), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n793), .A2(G317), .B1(new_n825), .B2(G303), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n766), .A2(G322), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n796), .C2(new_n774), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT49), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n768), .A2(new_n512), .B1(new_n777), .B2(new_n790), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n424), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1056), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1048), .B1(new_n1067), .B2(new_n763), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1034), .A2(new_n749), .B1(new_n1037), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1036), .A2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n995), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n989), .B(KEYINPUT44), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n684), .B1(new_n1072), .B2(new_n987), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n749), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n255), .A2(new_n805), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n803), .B1(new_n233), .B2(new_n519), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n750), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n791), .A2(new_n831), .B1(new_n396), .B2(new_n783), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT51), .Z(new_n1080));
  NOR2_X1   g0880(.A1(new_n798), .A2(new_n216), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G50), .B2(new_n773), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n210), .B2(new_n780), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n349), .A2(new_n825), .B1(new_n794), .B2(G143), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n424), .A3(new_n827), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1080), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT109), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G317), .A2(new_n766), .B1(new_n793), .B2(G311), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n257), .B1(new_n794), .B2(G322), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n497), .B2(new_n782), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n774), .A2(new_n532), .B1(new_n768), .B2(new_n218), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n798), .A2(new_n512), .B1(new_n780), .B2(new_n799), .ZN(new_n1094));
  OR4_X1    g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1088), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1078), .B1(new_n1097), .B2(new_n763), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n982), .B2(new_n759), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n691), .B1(new_n1035), .B2(new_n996), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1074), .B1(new_n744), .B2(new_n1034), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1075), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(KEYINPUT112), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n893), .A2(new_n895), .ZN(new_n1104));
  OAI211_X1 g0904(.A(KEYINPUT111), .B(G330), .C1(new_n929), .C2(new_n931), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n817), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT111), .B1(new_n939), .B2(G330), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1104), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n896), .A2(new_n742), .A3(G330), .A4(new_n817), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n816), .A2(new_n368), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n815), .B1(new_n699), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(G330), .B1(new_n929), .B2(new_n931), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT111), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n817), .A3(new_n1105), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1103), .B1(new_n1117), .B2(new_n1104), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT113), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT112), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT113), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1108), .A4(new_n1112), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1114), .A2(new_n933), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n817), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1104), .B1(new_n743), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n888), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT114), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n458), .A2(G330), .A3(new_n939), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n922), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1129), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1137), .B2(new_n1134), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n916), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n888), .B2(new_n1104), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n909), .A2(new_n1140), .A3(new_n912), .A4(new_n914), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n924), .B(new_n1139), .C1(new_n1111), .C2(new_n1104), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1125), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT110), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1109), .A3(new_n1142), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT110), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1147), .A3(new_n1125), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1136), .A2(new_n1138), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1147), .B1(new_n1143), .B2(new_n1125), .ZN(new_n1151));
  AOI211_X1 g0951(.A(KEYINPUT110), .B(new_n1126), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1146), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1134), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n692), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n915), .A2(new_n757), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n774), .A2(new_n830), .B1(new_n768), .B2(new_n202), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n791), .A2(new_n1160), .B1(new_n396), .B2(new_n798), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n783), .A2(new_n836), .B1(new_n782), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n625), .B(new_n1164), .C1(G125), .C2(new_n794), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1053), .A2(new_n780), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT53), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n766), .A2(G283), .B1(new_n825), .B2(new_n559), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n218), .B2(new_n774), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT115), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n625), .B1(new_n777), .B2(new_n497), .C1(new_n783), .C2(new_n512), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n210), .A2(new_n768), .B1(new_n780), .B2(new_n212), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n1172), .A2(new_n1081), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1168), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1175), .A2(new_n763), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n751), .B(new_n1176), .C1(new_n284), .C2(new_n844), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1158), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1149), .B2(new_n748), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1157), .A2(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n346), .A2(new_n299), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n342), .A2(new_n669), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G330), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n937), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1184), .B(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(G330), .C1(new_n940), .C2(new_n942), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(new_n919), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1186), .A2(new_n843), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n768), .A2(new_n283), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G97), .B2(new_n773), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n512), .B2(new_n791), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n793), .A2(G107), .B1(new_n825), .B2(new_n352), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n799), .B2(new_n777), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n804), .A2(new_n480), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n798), .A2(new_n210), .B1(new_n780), .B2(new_n216), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT118), .Z(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G33), .A2(G41), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT116), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n202), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT117), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n793), .A2(G128), .B1(new_n825), .B2(G137), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n780), .B2(new_n1163), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n798), .A2(new_n831), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n766), .A2(G125), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n774), .B2(new_n836), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1206), .B1(G124), .B2(new_n794), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1217), .B1(new_n396), .B2(new_n768), .C1(new_n1214), .C2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1204), .B(new_n1208), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n763), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT119), .Z(new_n1223));
  AOI211_X1 g1023(.A(new_n751), .B(new_n1223), .C1(new_n202), .C2(new_n844), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1193), .A2(new_n749), .B1(new_n1194), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1135), .B1(new_n1149), .B2(new_n1137), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(KEYINPUT57), .A3(new_n1193), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n691), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1193), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1137), .A2(new_n1134), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1005), .B(KEYINPUT120), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1136), .A2(new_n1138), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n896), .A2(new_n757), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n512), .A2(new_n774), .B1(new_n791), .B2(new_n497), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G97), .B2(new_n822), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1049), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n783), .A2(new_n799), .B1(new_n782), .B2(new_n218), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n257), .B(new_n1238), .C1(G303), .C2(new_n794), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n961), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n822), .A2(G159), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n202), .B2(new_n798), .C1(new_n774), .C2(new_n1163), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n782), .A2(new_n831), .B1(new_n777), .B2(new_n1160), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G137), .B2(new_n793), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1195), .B1(G132), .B2(new_n766), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n424), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n763), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n751), .B1(new_n844), .B2(new_n210), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1137), .A2(new_n748), .B1(new_n1234), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1233), .A2(new_n1252), .ZN(G381));
  AOI21_X1  g1053(.A(new_n1030), .B1(new_n1074), .B2(new_n1034), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n748), .B1(new_n1254), .B2(new_n1005), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1027), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n1025), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1255), .A2(new_n1257), .B1(new_n956), .B2(new_n977), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1075), .A2(new_n1099), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1100), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1101), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G396), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1036), .A2(new_n1263), .A3(new_n1069), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1258), .A2(new_n847), .A3(new_n1262), .A4(new_n1265), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1266), .ZN(G407));
  AOI21_X1  g1067(.A(new_n1179), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n670), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(G375), .C2(new_n1271), .ZN(G409));
  INV_X1    g1072(.A(KEYINPUT123), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1258), .B2(G390), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1263), .B1(new_n1036), .B2(new_n1069), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1265), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(G387), .A2(new_n1262), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n1278), .B2(new_n978), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1274), .A2(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1258), .A2(G390), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1262), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1265), .A2(new_n1275), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1273), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1226), .A2(new_n1193), .A3(new_n1232), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1225), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1268), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT121), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1225), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(KEYINPUT121), .A3(new_n1268), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1124), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1134), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n691), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1134), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1231), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n847), .B1(new_n1298), .B2(new_n1251), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1297), .A2(new_n1231), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G384), .B(new_n1252), .C1(new_n1300), .C2(new_n1296), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1293), .A2(new_n1294), .A3(new_n1269), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1287), .A2(KEYINPUT121), .A3(new_n1268), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT121), .B1(new_n1287), .B2(new_n1268), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1270), .B1(new_n1308), .B2(new_n1291), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1270), .A2(KEYINPUT122), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1299), .A2(new_n1301), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1270), .A2(G2897), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1311), .B(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1304), .B(new_n1305), .C1(new_n1309), .C2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1294), .B1(new_n1309), .B2(new_n1303), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1285), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1309), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1303), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1293), .A2(new_n1269), .A3(new_n1303), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1280), .A2(new_n1305), .A3(new_n1284), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(KEYINPUT124), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1293), .A2(new_n1269), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1311), .B(new_n1312), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1318), .A2(new_n1322), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1317), .A2(new_n1329), .ZN(G405));
  INV_X1    g1130(.A(KEYINPUT57), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1134), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1332));
  XOR2_X1   g1132(.A(new_n1192), .B(new_n919), .Z(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(new_n691), .A3(new_n1227), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1335), .A2(G378), .A3(new_n1225), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G378), .B1(new_n1335), .B2(new_n1225), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1303), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT126), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(KEYINPUT126), .B(new_n1303), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G375), .A2(new_n1268), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1343), .A2(new_n1291), .A3(new_n1302), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1343), .A2(KEYINPUT127), .A3(new_n1291), .A4(new_n1302), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1342), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1285), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1342), .A2(new_n1348), .A3(new_n1284), .A4(new_n1280), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


