

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771;

  NOR2_X2 U371 ( .A1(n688), .A2(n687), .ZN(n651) );
  XNOR2_X1 U372 ( .A(n580), .B(KEYINPUT105), .ZN(n764) );
  AND2_X1 U373 ( .A1(n388), .A2(n398), .ZN(n353) );
  XNOR2_X1 U374 ( .A(n608), .B(KEYINPUT100), .ZN(n680) );
  XNOR2_X1 U375 ( .A(n475), .B(n474), .ZN(n552) );
  XOR2_X1 U376 ( .A(G113), .B(G104), .Z(n561) );
  XNOR2_X1 U377 ( .A(n489), .B(G122), .ZN(n556) );
  INV_X1 U378 ( .A(G107), .ZN(n489) );
  AND2_X2 U379 ( .A1(n402), .A2(n459), .ZN(n454) );
  XNOR2_X1 U380 ( .A(n478), .B(n558), .ZN(n477) );
  AND2_X2 U381 ( .A1(n740), .A2(n366), .ZN(n464) );
  INV_X2 U382 ( .A(G953), .ZN(n755) );
  XNOR2_X2 U383 ( .A(n397), .B(n522), .ZN(n659) );
  BUF_X1 U384 ( .A(n587), .Z(n614) );
  XNOR2_X1 U385 ( .A(n454), .B(KEYINPUT48), .ZN(n453) );
  NOR2_X1 U386 ( .A1(n767), .A2(n452), .ZN(n451) );
  INV_X1 U387 ( .A(n686), .ZN(n452) );
  NOR2_X1 U388 ( .A1(n581), .A2(n380), .ZN(n582) );
  NOR2_X1 U389 ( .A1(n587), .A2(n484), .ZN(n483) );
  INV_X1 U390 ( .A(G131), .ZN(n495) );
  XOR2_X1 U391 ( .A(KEYINPUT4), .B(G146), .Z(n537) );
  AND2_X1 U392 ( .A1(n408), .A2(n365), .ZN(n433) );
  AND2_X2 U393 ( .A1(n453), .A2(n451), .ZN(n753) );
  AND2_X1 U394 ( .A1(n377), .A2(n376), .ZN(n375) );
  OR2_X1 U395 ( .A1(n620), .A2(n372), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n483), .B(KEYINPUT19), .ZN(n620) );
  XNOR2_X1 U397 ( .A(n560), .B(n559), .ZN(n606) );
  OR2_X1 U398 ( .A1(n661), .A2(G902), .ZN(n407) );
  XNOR2_X1 U399 ( .A(n537), .B(n494), .ZN(n493) );
  XNOR2_X1 U400 ( .A(n487), .B(G110), .ZN(n531) );
  XNOR2_X1 U401 ( .A(n495), .B(G137), .ZN(n494) );
  BUF_X1 U402 ( .A(n368), .Z(n349) );
  BUF_X1 U403 ( .A(n731), .Z(n350) );
  NAND2_X1 U404 ( .A1(n390), .A2(n433), .ZN(n351) );
  NAND2_X1 U405 ( .A1(n390), .A2(n433), .ZN(n432) );
  XNOR2_X1 U406 ( .A(n556), .B(n534), .ZN(n488) );
  XNOR2_X1 U407 ( .A(KEYINPUT16), .B(KEYINPUT70), .ZN(n534) );
  NAND2_X1 U408 ( .A1(n482), .A2(n492), .ZN(n391) );
  INV_X1 U409 ( .A(G472), .ZN(n381) );
  INV_X1 U410 ( .A(n694), .ZN(n429) );
  INV_X1 U411 ( .A(KEYINPUT8), .ZN(n474) );
  NAND2_X1 U412 ( .A1(n755), .A2(G234), .ZN(n475) );
  OR2_X2 U413 ( .A1(n753), .A2(KEYINPUT78), .ZN(n408) );
  INV_X1 U414 ( .A(KEYINPUT72), .ZN(n389) );
  XNOR2_X1 U415 ( .A(n533), .B(n485), .ZN(n736) );
  XNOR2_X1 U416 ( .A(n488), .B(n486), .ZN(n485) );
  INV_X1 U417 ( .A(n531), .ZN(n486) );
  NOR2_X1 U418 ( .A1(n384), .A2(n383), .ZN(n421) );
  INV_X1 U419 ( .A(G134), .ZN(n496) );
  AND2_X1 U420 ( .A1(n399), .A2(n680), .ZN(n398) );
  INV_X1 U421 ( .A(n581), .ZN(n399) );
  NAND2_X1 U422 ( .A1(n530), .A2(n472), .ZN(n470) );
  NOR2_X1 U423 ( .A1(n626), .A2(n631), .ZN(n435) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n434) );
  INV_X1 U425 ( .A(KEYINPUT22), .ZN(n624) );
  XOR2_X1 U426 ( .A(n646), .B(KEYINPUT101), .Z(n530) );
  XNOR2_X1 U427 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U428 ( .A(KEYINPUT30), .ZN(n410) );
  XNOR2_X1 U429 ( .A(n574), .B(n406), .ZN(n405) );
  INV_X1 U430 ( .A(G475), .ZN(n406) );
  NOR2_X1 U431 ( .A1(n729), .A2(G902), .ZN(n560) );
  XNOR2_X1 U432 ( .A(n614), .B(n458), .ZN(n473) );
  INV_X1 U433 ( .A(KEYINPUT38), .ZN(n458) );
  XNOR2_X1 U434 ( .A(G143), .B(G131), .ZN(n562) );
  XNOR2_X1 U435 ( .A(G122), .B(KEYINPUT93), .ZN(n563) );
  XOR2_X1 U436 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n564) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(KEYINPUT11), .Z(n569) );
  NAND2_X1 U438 ( .A1(G902), .A2(G469), .ZN(n417) );
  NAND2_X1 U439 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U440 ( .A(G469), .ZN(n415) );
  INV_X1 U441 ( .A(G902), .ZN(n414) );
  XNOR2_X1 U442 ( .A(KEYINPUT5), .B(KEYINPUT89), .ZN(n523) );
  XNOR2_X1 U443 ( .A(KEYINPUT88), .B(KEYINPUT73), .ZN(n524) );
  XOR2_X1 U444 ( .A(G113), .B(G119), .Z(n525) );
  NOR2_X1 U445 ( .A1(G953), .A2(G237), .ZN(n567) );
  AND2_X1 U446 ( .A1(n611), .A2(n357), .ZN(n402) );
  XOR2_X1 U447 ( .A(KEYINPUT3), .B(G116), .Z(n532) );
  NOR2_X1 U448 ( .A1(n694), .A2(KEYINPUT99), .ZN(n422) );
  XNOR2_X1 U449 ( .A(G125), .B(KEYINPUT82), .ZN(n535) );
  XOR2_X1 U450 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n536) );
  INV_X1 U451 ( .A(KEYINPUT83), .ZN(n541) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n499) );
  OR2_X1 U453 ( .A1(G237), .A2(G902), .ZN(n548) );
  INV_X1 U454 ( .A(n473), .ZN(n472) );
  OR2_X1 U455 ( .A1(n352), .A2(n551), .ZN(n467) );
  XNOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n497) );
  XNOR2_X1 U457 ( .A(n513), .B(KEYINPUT25), .ZN(n490) );
  OR2_X1 U458 ( .A1(n733), .A2(G902), .ZN(n491) );
  NOR2_X1 U459 ( .A1(n703), .A2(n702), .ZN(n699) );
  XOR2_X1 U460 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n508) );
  INV_X1 U461 ( .A(G119), .ZN(n487) );
  XNOR2_X1 U462 ( .A(G107), .B(G110), .ZN(n516) );
  XOR2_X1 U463 ( .A(G140), .B(KEYINPUT87), .Z(n517) );
  INV_X1 U464 ( .A(KEYINPUT90), .ZN(n385) );
  NOR2_X1 U465 ( .A1(n630), .A2(n449), .ZN(n642) );
  XNOR2_X1 U466 ( .A(n555), .B(n477), .ZN(n729) );
  XOR2_X1 U467 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n554) );
  INV_X1 U468 ( .A(KEYINPUT42), .ZN(n455) );
  XNOR2_X1 U469 ( .A(n610), .B(n462), .ZN(n769) );
  NAND2_X1 U470 ( .A1(n476), .A2(n449), .ZN(n580) );
  XNOR2_X1 U471 ( .A(n404), .B(n579), .ZN(n476) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n393) );
  INV_X1 U473 ( .A(n636), .ZN(n395) );
  INV_X1 U474 ( .A(KEYINPUT32), .ZN(n628) );
  NAND2_X1 U475 ( .A1(n352), .A2(n530), .ZN(n593) );
  INV_X1 U476 ( .A(KEYINPUT56), .ZN(n439) );
  AND2_X1 U477 ( .A1(n409), .A2(n577), .ZN(n352) );
  NAND2_X1 U478 ( .A1(n642), .A2(n378), .ZN(n427) );
  INV_X1 U479 ( .A(n427), .ZN(n425) );
  XOR2_X1 U480 ( .A(G902), .B(KEYINPUT15), .Z(n547) );
  XOR2_X1 U481 ( .A(n544), .B(n543), .Z(n354) );
  XOR2_X1 U482 ( .A(n529), .B(n528), .Z(n355) );
  XOR2_X1 U483 ( .A(G137), .B(G128), .Z(n356) );
  AND2_X1 U484 ( .A1(n591), .A2(n590), .ZN(n357) );
  NOR2_X1 U485 ( .A1(n710), .A2(n387), .ZN(n358) );
  AND2_X1 U486 ( .A1(n472), .A2(n471), .ZN(n359) );
  OR2_X1 U487 ( .A1(n427), .A2(KEYINPUT99), .ZN(n360) );
  XOR2_X1 U488 ( .A(n726), .B(n725), .Z(n361) );
  XOR2_X1 U489 ( .A(n663), .B(n662), .Z(n362) );
  XNOR2_X1 U490 ( .A(n659), .B(n658), .ZN(n363) );
  XOR2_X1 U491 ( .A(n654), .B(n653), .Z(n364) );
  INV_X1 U492 ( .A(KEYINPUT99), .ZN(n437) );
  INV_X1 U493 ( .A(KEYINPUT78), .ZN(n492) );
  OR2_X1 U494 ( .A1(n650), .A2(n687), .ZN(n365) );
  AND2_X1 U495 ( .A1(n547), .A2(KEYINPUT78), .ZN(n366) );
  INV_X1 U496 ( .A(n735), .ZN(n444) );
  XOR2_X1 U497 ( .A(n665), .B(KEYINPUT60), .Z(n367) );
  AND2_X2 U498 ( .A1(n432), .A2(n431), .ZN(n368) );
  AND2_X2 U499 ( .A1(n351), .A2(n431), .ZN(n731) );
  NAND2_X1 U500 ( .A1(n375), .A2(n374), .ZN(n369) );
  NAND2_X1 U501 ( .A1(n375), .A2(n374), .ZN(n643) );
  XNOR2_X1 U502 ( .A(n549), .B(n498), .ZN(n587) );
  XNOR2_X1 U503 ( .A(n481), .B(n633), .ZN(n638) );
  OR2_X1 U504 ( .A1(n412), .A2(n416), .ZN(n370) );
  AND2_X1 U505 ( .A1(n473), .A2(n484), .ZN(n691) );
  OR2_X2 U506 ( .A1(n607), .A2(n717), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(KEYINPUT41), .ZN(n717) );
  OR2_X1 U508 ( .A1(n473), .A2(n484), .ZN(n604) );
  INV_X1 U509 ( .A(n677), .ZN(n371) );
  NAND2_X1 U510 ( .A1(n419), .A2(n421), .ZN(n649) );
  NAND2_X1 U511 ( .A1(n420), .A2(n637), .ZN(n419) );
  XNOR2_X1 U512 ( .A(n480), .B(KEYINPUT44), .ZN(n420) );
  OR2_X2 U513 ( .A1(n416), .A2(n412), .ZN(n583) );
  XNOR2_X1 U514 ( .A(n511), .B(n573), .ZN(n733) );
  XNOR2_X1 U515 ( .A(n634), .B(n389), .ZN(n382) );
  OR2_X1 U516 ( .A1(n619), .A2(KEYINPUT0), .ZN(n372) );
  AND2_X1 U517 ( .A1(n641), .A2(n631), .ZN(n378) );
  INV_X1 U518 ( .A(n641), .ZN(n388) );
  BUF_X1 U519 ( .A(n708), .Z(n379) );
  XNOR2_X1 U520 ( .A(n708), .B(KEYINPUT6), .ZN(n641) );
  XNOR2_X1 U521 ( .A(n583), .B(n497), .ZN(n373) );
  XNOR2_X1 U522 ( .A(n583), .B(n497), .ZN(n698) );
  NOR2_X1 U523 ( .A1(n643), .A2(n623), .ZN(n625) );
  NAND2_X1 U524 ( .A1(n619), .A2(KEYINPUT0), .ZN(n376) );
  NAND2_X1 U525 ( .A1(n620), .A2(KEYINPUT0), .ZN(n377) );
  NAND2_X1 U526 ( .A1(n708), .A2(n690), .ZN(n411) );
  INV_X1 U527 ( .A(n708), .ZN(n380) );
  XNOR2_X2 U528 ( .A(n463), .B(n381), .ZN(n708) );
  AND2_X2 U529 ( .A1(n382), .A2(n388), .ZN(n448) );
  NAND2_X1 U530 ( .A1(n382), .A2(n379), .ZN(n386) );
  NAND2_X1 U531 ( .A1(n768), .A2(n673), .ZN(n481) );
  NAND2_X1 U532 ( .A1(n640), .A2(n426), .ZN(n383) );
  NAND2_X1 U533 ( .A1(n423), .A2(n360), .ZN(n384) );
  XNOR2_X2 U534 ( .A(n386), .B(n385), .ZN(n387) );
  NAND2_X1 U535 ( .A1(n430), .A2(n429), .ZN(n428) );
  XNOR2_X1 U536 ( .A(n648), .B(KEYINPUT91), .ZN(n430) );
  NAND2_X1 U537 ( .A1(n387), .A2(n645), .ZN(n644) );
  AND2_X2 U538 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U539 ( .A1(n464), .A2(n753), .ZN(n392) );
  NAND2_X1 U540 ( .A1(n763), .A2(n638), .ZN(n480) );
  XNOR2_X2 U541 ( .A(n394), .B(n393), .ZN(n763) );
  NAND2_X1 U542 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U543 ( .A(n635), .B(KEYINPUT34), .ZN(n396) );
  XNOR2_X1 U544 ( .A(n397), .B(n355), .ZN(n652) );
  XNOR2_X2 U545 ( .A(n752), .B(n538), .ZN(n397) );
  NAND2_X1 U546 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U547 ( .A(n764), .B(KEYINPUT79), .ZN(n591) );
  NAND2_X1 U548 ( .A1(n400), .A2(KEYINPUT65), .ZN(n640) );
  NAND2_X1 U549 ( .A1(n639), .A2(KEYINPUT44), .ZN(n400) );
  NOR2_X2 U550 ( .A1(n630), .A2(n627), .ZN(n629) );
  XNOR2_X1 U551 ( .A(n736), .B(n546), .ZN(n450) );
  NAND2_X1 U552 ( .A1(n401), .A2(n436), .ZN(n461) );
  INV_X1 U553 ( .A(n770), .ZN(n401) );
  XNOR2_X2 U554 ( .A(n456), .B(n455), .ZN(n770) );
  NAND2_X1 U555 ( .A1(n353), .A2(n690), .ZN(n612) );
  NAND2_X1 U556 ( .A1(n353), .A2(n403), .ZN(n404) );
  NOR2_X1 U557 ( .A1(n614), .A2(n484), .ZN(n403) );
  XNOR2_X2 U558 ( .A(n407), .B(n405), .ZN(n592) );
  XNOR2_X1 U559 ( .A(n572), .B(n573), .ZN(n661) );
  NOR2_X1 U560 ( .A1(n652), .A2(G902), .ZN(n463) );
  NOR2_X1 U561 ( .A1(n659), .A2(n413), .ZN(n412) );
  NAND2_X1 U562 ( .A1(n659), .A2(G469), .ZN(n418) );
  NAND2_X1 U563 ( .A1(n430), .A2(n422), .ZN(n426) );
  NAND2_X1 U564 ( .A1(n428), .A2(n424), .ZN(n423) );
  NOR2_X1 U565 ( .A1(n425), .A2(n437), .ZN(n424) );
  INV_X1 U566 ( .A(n651), .ZN(n431) );
  XNOR2_X1 U567 ( .A(n435), .B(n434), .ZN(n627) );
  NAND2_X1 U568 ( .A1(n552), .A2(G221), .ZN(n507) );
  INV_X1 U569 ( .A(n769), .ZN(n436) );
  XNOR2_X1 U570 ( .A(n438), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U571 ( .A1(n443), .A2(n444), .ZN(n438) );
  XNOR2_X1 U572 ( .A(n440), .B(n439), .ZN(G51) );
  NAND2_X1 U573 ( .A1(n447), .A2(n444), .ZN(n440) );
  XNOR2_X1 U574 ( .A(n441), .B(n367), .ZN(G60) );
  NAND2_X1 U575 ( .A1(n446), .A2(n444), .ZN(n441) );
  XNOR2_X1 U576 ( .A(n442), .B(KEYINPUT119), .ZN(G54) );
  NAND2_X1 U577 ( .A1(n445), .A2(n444), .ZN(n442) );
  XNOR2_X1 U578 ( .A(n655), .B(n364), .ZN(n443) );
  NAND2_X1 U579 ( .A1(n731), .A2(G472), .ZN(n655) );
  XNOR2_X1 U580 ( .A(n660), .B(n363), .ZN(n445) );
  XNOR2_X1 U581 ( .A(n664), .B(n362), .ZN(n446) );
  XNOR2_X1 U582 ( .A(n727), .B(n361), .ZN(n447) );
  XNOR2_X2 U583 ( .A(n448), .B(KEYINPUT33), .ZN(n718) );
  NOR2_X2 U584 ( .A1(n683), .A2(n670), .ZN(n648) );
  BUF_X2 U585 ( .A(n373), .Z(n449) );
  NOR2_X1 U586 ( .A1(n450), .A2(n547), .ZN(n549) );
  XNOR2_X1 U587 ( .A(n450), .B(KEYINPUT55), .ZN(n725) );
  NOR2_X1 U588 ( .A1(n693), .A2(n692), .ZN(n457) );
  XNOR2_X1 U589 ( .A(n461), .B(n460), .ZN(n459) );
  INV_X1 U590 ( .A(KEYINPUT46), .ZN(n460) );
  INV_X1 U591 ( .A(KEYINPUT40), .ZN(n462) );
  NAND2_X1 U592 ( .A1(n466), .A2(n465), .ZN(n609) );
  NAND2_X1 U593 ( .A1(n470), .A2(n551), .ZN(n465) );
  NAND2_X1 U594 ( .A1(n468), .A2(n467), .ZN(n466) );
  NAND2_X1 U595 ( .A1(n352), .A2(n469), .ZN(n468) );
  NAND2_X1 U596 ( .A1(n359), .A2(n530), .ZN(n469) );
  INV_X1 U597 ( .A(n551), .ZN(n471) );
  NAND2_X1 U598 ( .A1(n552), .A2(G217), .ZN(n553) );
  XNOR2_X1 U599 ( .A(n557), .B(n479), .ZN(n478) );
  INV_X1 U600 ( .A(KEYINPUT96), .ZN(n479) );
  NOR2_X2 U601 ( .A1(n606), .A2(n592), .ZN(n608) );
  NAND2_X1 U602 ( .A1(n740), .A2(n547), .ZN(n482) );
  XNOR2_X2 U603 ( .A(n649), .B(KEYINPUT45), .ZN(n740) );
  INV_X1 U604 ( .A(n614), .ZN(n595) );
  INV_X1 U605 ( .A(n690), .ZN(n484) );
  XNOR2_X2 U606 ( .A(n491), .B(n490), .ZN(n703) );
  NAND2_X1 U607 ( .A1(n740), .A2(n753), .ZN(n688) );
  XNOR2_X2 U608 ( .A(n558), .B(n493), .ZN(n752) );
  XNOR2_X2 U609 ( .A(n544), .B(n496), .ZN(n558) );
  XNOR2_X2 U610 ( .A(n521), .B(G128), .ZN(n544) );
  NAND2_X1 U611 ( .A1(n698), .A2(n699), .ZN(n634) );
  AND2_X1 U612 ( .A1(G210), .A2(n548), .ZN(n498) );
  XNOR2_X1 U613 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n545), .B(n354), .ZN(n546) );
  INV_X1 U615 ( .A(n702), .ZN(n621) );
  NAND2_X1 U616 ( .A1(n622), .A2(n621), .ZN(n623) );
  INV_X1 U617 ( .A(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT39), .ZN(n551) );
  INV_X1 U619 ( .A(KEYINPUT121), .ZN(n665) );
  NOR2_X1 U620 ( .A1(G952), .A2(n755), .ZN(n735) );
  XNOR2_X1 U621 ( .A(n499), .B(KEYINPUT14), .ZN(n501) );
  NAND2_X1 U622 ( .A1(n501), .A2(G952), .ZN(n500) );
  XNOR2_X1 U623 ( .A(n500), .B(KEYINPUT84), .ZN(n716) );
  NOR2_X1 U624 ( .A1(G953), .A2(n716), .ZN(n618) );
  NAND2_X1 U625 ( .A1(n501), .A2(G902), .ZN(n502) );
  XNOR2_X1 U626 ( .A(KEYINPUT86), .B(n502), .ZN(n616) );
  OR2_X1 U627 ( .A1(n616), .A2(n755), .ZN(n503) );
  NOR2_X1 U628 ( .A1(G900), .A2(n503), .ZN(n504) );
  NOR2_X1 U629 ( .A1(n618), .A2(n504), .ZN(n505) );
  XNOR2_X1 U630 ( .A(KEYINPUT75), .B(n505), .ZN(n577) );
  XOR2_X1 U631 ( .A(G125), .B(G140), .Z(n506) );
  XNOR2_X1 U632 ( .A(KEYINPUT10), .B(n506), .ZN(n751) );
  XNOR2_X1 U633 ( .A(G146), .B(n751), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U635 ( .A(n531), .B(n356), .ZN(n509) );
  XNOR2_X1 U636 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U637 ( .A(n547), .ZN(n650) );
  NAND2_X1 U638 ( .A1(n650), .A2(G234), .ZN(n512) );
  XNOR2_X1 U639 ( .A(n512), .B(KEYINPUT20), .ZN(n514) );
  NAND2_X1 U640 ( .A1(G217), .A2(n514), .ZN(n513) );
  NAND2_X1 U641 ( .A1(G221), .A2(n514), .ZN(n515) );
  XNOR2_X1 U642 ( .A(KEYINPUT21), .B(n515), .ZN(n702) );
  XNOR2_X1 U643 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U644 ( .A(G104), .B(n518), .Z(n520) );
  NAND2_X1 U645 ( .A1(G227), .A2(n755), .ZN(n519) );
  XNOR2_X1 U646 ( .A(n520), .B(n519), .ZN(n522) );
  XNOR2_X2 U647 ( .A(G143), .B(KEYINPUT64), .ZN(n521) );
  XOR2_X2 U648 ( .A(KEYINPUT68), .B(G101), .Z(n538) );
  AND2_X1 U649 ( .A1(n370), .A2(n699), .ZN(n646) );
  NAND2_X1 U650 ( .A1(G214), .A2(n548), .ZN(n690) );
  XNOR2_X1 U651 ( .A(n523), .B(n532), .ZN(n527) );
  XNOR2_X1 U652 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U653 ( .A(n527), .B(n526), .Z(n529) );
  NAND2_X1 U654 ( .A1(n567), .A2(G210), .ZN(n528) );
  XNOR2_X1 U655 ( .A(n532), .B(n561), .ZN(n533) );
  XOR2_X1 U656 ( .A(n536), .B(n535), .Z(n540) );
  XNOR2_X1 U657 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U658 ( .A(n540), .B(n539), .ZN(n545) );
  NAND2_X1 U659 ( .A1(G224), .A2(n755), .ZN(n542) );
  INV_X1 U660 ( .A(KEYINPUT69), .ZN(n550) );
  XNOR2_X1 U661 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U662 ( .A(n556), .B(G116), .ZN(n557) );
  XNOR2_X1 U663 ( .A(KEYINPUT97), .B(G478), .ZN(n559) );
  XNOR2_X1 U664 ( .A(n562), .B(n561), .ZN(n566) );
  XNOR2_X1 U665 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U666 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U667 ( .A1(G214), .A2(n567), .ZN(n568) );
  XNOR2_X1 U668 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U669 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U670 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n606), .A2(n592), .ZN(n575) );
  XOR2_X1 U672 ( .A(KEYINPUT98), .B(n575), .Z(n682) );
  AND2_X1 U673 ( .A1(n609), .A2(n682), .ZN(n576) );
  XNOR2_X1 U674 ( .A(n576), .B(KEYINPUT106), .ZN(n767) );
  XNOR2_X1 U675 ( .A(KEYINPUT81), .B(KEYINPUT36), .ZN(n579) );
  INV_X1 U676 ( .A(n703), .ZN(n631) );
  NOR2_X1 U677 ( .A1(n702), .A2(n631), .ZN(n578) );
  NAND2_X1 U678 ( .A1(n578), .A2(n577), .ZN(n581) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(n582), .ZN(n585) );
  XNOR2_X1 U680 ( .A(n370), .B(KEYINPUT102), .ZN(n584) );
  NAND2_X1 U681 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U682 ( .A(KEYINPUT103), .B(n586), .Z(n607) );
  NOR2_X1 U683 ( .A1(n607), .A2(n620), .ZN(n677) );
  INV_X1 U684 ( .A(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n677), .A2(n588), .ZN(n589) );
  NAND2_X1 U686 ( .A1(KEYINPUT47), .A2(n589), .ZN(n590) );
  INV_X1 U687 ( .A(n592), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n636) );
  NOR2_X1 U689 ( .A1(n593), .A2(n636), .ZN(n594) );
  NAND2_X1 U690 ( .A1(n595), .A2(n594), .ZN(n676) );
  NOR2_X1 U691 ( .A1(n608), .A2(n682), .ZN(n694) );
  NAND2_X1 U692 ( .A1(KEYINPUT47), .A2(n694), .ZN(n596) );
  XOR2_X1 U693 ( .A(KEYINPUT77), .B(n596), .Z(n597) );
  NAND2_X1 U694 ( .A1(n676), .A2(n597), .ZN(n598) );
  XNOR2_X1 U695 ( .A(n598), .B(KEYINPUT76), .ZN(n603) );
  XNOR2_X1 U696 ( .A(KEYINPUT71), .B(n694), .ZN(n600) );
  INV_X1 U697 ( .A(KEYINPUT47), .ZN(n599) );
  NAND2_X1 U698 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U699 ( .A1(n371), .A2(n601), .ZN(n602) );
  NOR2_X1 U700 ( .A1(n603), .A2(n602), .ZN(n611) );
  XNOR2_X1 U701 ( .A(KEYINPUT104), .B(n604), .ZN(n693) );
  NOR2_X1 U702 ( .A1(n606), .A2(n605), .ZN(n622) );
  INV_X1 U703 ( .A(n622), .ZN(n692) );
  NAND2_X1 U704 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U705 ( .A1(n612), .A2(n449), .ZN(n613) );
  XNOR2_X1 U706 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  NAND2_X1 U707 ( .A1(n615), .A2(n614), .ZN(n686) );
  INV_X1 U708 ( .A(KEYINPUT80), .ZN(n633) );
  XNOR2_X1 U709 ( .A(G898), .B(KEYINPUT85), .ZN(n743) );
  NAND2_X1 U710 ( .A1(G953), .A2(n743), .ZN(n738) );
  NOR2_X1 U711 ( .A1(n616), .A2(n738), .ZN(n617) );
  NOR2_X1 U712 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U713 ( .A(n625), .B(n624), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n449), .A2(n641), .ZN(n626) );
  XNOR2_X2 U715 ( .A(n629), .B(n628), .ZN(n768) );
  NOR2_X1 U716 ( .A1(n379), .A2(n631), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n642), .A2(n632), .ZN(n673) );
  NOR2_X1 U718 ( .A1(n369), .A2(n718), .ZN(n635) );
  NAND2_X1 U719 ( .A1(KEYINPUT65), .A2(n763), .ZN(n637) );
  INV_X1 U720 ( .A(n638), .ZN(n639) );
  INV_X1 U721 ( .A(n369), .ZN(n645) );
  XNOR2_X2 U722 ( .A(n644), .B(KEYINPUT31), .ZN(n683) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n379), .A2(n647), .ZN(n670) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n687) );
  XNOR2_X1 U726 ( .A(n652), .B(KEYINPUT107), .ZN(n654) );
  XOR2_X1 U727 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n368), .A2(G469), .ZN(n660) );
  XNOR2_X1 U731 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n661), .B(KEYINPUT120), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n368), .A2(G475), .ZN(n664) );
  XOR2_X1 U734 ( .A(G101), .B(n425), .Z(G3) );
  NAND2_X1 U735 ( .A1(n680), .A2(n670), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(G104), .ZN(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n668) );
  XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT108), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U740 ( .A(KEYINPUT26), .B(n669), .Z(n672) );
  NAND2_X1 U741 ( .A1(n670), .A2(n682), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G9) );
  XNOR2_X1 U743 ( .A(G110), .B(n673), .ZN(G12) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U745 ( .A1(n677), .A2(n682), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(G30) );
  XNOR2_X1 U747 ( .A(G143), .B(n676), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n680), .A2(n677), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n678), .B(KEYINPUT110), .ZN(n679) );
  XNOR2_X1 U750 ( .A(G146), .B(n679), .ZN(G48) );
  NAND2_X1 U751 ( .A1(n680), .A2(n683), .ZN(n681) );
  XNOR2_X1 U752 ( .A(n681), .B(G113), .ZN(G15) );
  XOR2_X1 U753 ( .A(G116), .B(KEYINPUT111), .Z(n685) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(G18) );
  XNOR2_X1 U756 ( .A(G140), .B(n686), .ZN(G42) );
  XNOR2_X1 U757 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n689), .A2(n755), .ZN(n723) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U762 ( .A1(n718), .A2(n697), .ZN(n713) );
  XNOR2_X1 U763 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n699), .A2(n449), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n701), .B(n700), .ZN(n706) );
  NAND2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n704), .Z(n705) );
  NAND2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U770 ( .A(n709), .B(KEYINPUT114), .ZN(n710) );
  XOR2_X1 U771 ( .A(KEYINPUT51), .B(n358), .Z(n711) );
  NOR2_X1 U772 ( .A1(n717), .A2(n711), .ZN(n712) );
  NOR2_X1 U773 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U774 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT115), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U780 ( .A(KEYINPUT53), .B(n724), .ZN(G75) );
  XOR2_X1 U781 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n726) );
  NAND2_X1 U782 ( .A1(n731), .A2(G210), .ZN(n727) );
  NAND2_X1 U783 ( .A1(G478), .A2(n349), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n735), .A2(n730), .ZN(G63) );
  NAND2_X1 U786 ( .A1(G217), .A2(n350), .ZN(n732) );
  XNOR2_X1 U787 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U788 ( .A1(n735), .A2(n734), .ZN(G66) );
  XOR2_X1 U789 ( .A(n736), .B(KEYINPUT123), .Z(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(G101), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n750) );
  AND2_X1 U792 ( .A1(n740), .A2(n755), .ZN(n746) );
  XOR2_X1 U793 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n742) );
  NAND2_X1 U794 ( .A1(G224), .A2(G953), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n742), .B(n741), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U798 ( .A(n747), .B(KEYINPUT124), .Z(n748) );
  XNOR2_X1 U799 ( .A(KEYINPUT125), .B(n748), .ZN(n749) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U801 ( .A(n752), .B(n751), .Z(n757) );
  INV_X1 U802 ( .A(n757), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n762) );
  XNOR2_X1 U805 ( .A(G227), .B(KEYINPUT126), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G900), .A2(n759), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(G953), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U810 ( .A(n763), .B(G122), .ZN(G24) );
  XNOR2_X1 U811 ( .A(n764), .B(G125), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n765), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U813 ( .A(G134), .B(KEYINPUT112), .Z(n766) );
  XNOR2_X1 U814 ( .A(n767), .B(n766), .ZN(G36) );
  XNOR2_X1 U815 ( .A(n768), .B(G119), .ZN(G21) );
  XOR2_X1 U816 ( .A(G131), .B(n769), .Z(G33) );
  XNOR2_X1 U817 ( .A(G137), .B(KEYINPUT127), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n771), .B(n770), .ZN(G39) );
endmodule

