//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n551, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NAND3_X1  g047(.A1(new_n465), .A2(G124), .A3(G2105), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n464), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n464), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n473), .B(new_n475), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(new_n476), .A2(G138), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n464), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n460), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G102), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n486), .A2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT6), .A3(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AND4_X1   g076(.A1(new_n495), .A2(new_n501), .A3(G50), .A4(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n498), .B2(new_n500), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n495), .B1(new_n504), .B2(G50), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n498), .B2(new_n500), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n509), .A3(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G88), .B1(new_n514), .B2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n506), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n511), .A2(G89), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n504), .A2(G51), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  NAND2_X1  g100(.A1(G77), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n510), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT69), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n501), .A2(new_n520), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n501), .A2(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n510), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT72), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT73), .B(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n511), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n504), .A2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n533), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n504), .A2(KEYINPUT9), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n508), .A2(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT74), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(G65), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n497), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n511), .A2(G91), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n560), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n511), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n504), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AND2_X1   g151(.A1(new_n520), .A2(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT76), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n504), .A2(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n511), .A2(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G305));
  NAND3_X1  g158(.A1(new_n501), .A2(G85), .A3(new_n520), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n501), .A2(G47), .A3(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n497), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n510), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n593), .A2(KEYINPUT77), .A3(new_n584), .A4(new_n585), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n589), .A2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n511), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n564), .A2(G66), .A3(new_n565), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n504), .A2(G54), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT78), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n497), .B1(new_n601), .B2(new_n602), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n608));
  INV_X1    g183(.A(new_n605), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT79), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n597), .B1(new_n612), .B2(new_n596), .ZN(G284));
  AOI21_X1  g188(.A(new_n597), .B1(new_n612), .B2(new_n596), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n571), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n571), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n618), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n465), .A2(new_n491), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n465), .A2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G135), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n480), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2435), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2438), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(G14), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2100), .Z(new_n657));
  AND2_X1   g232(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT18), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n672), .B(new_n673), .C1(new_n671), .C2(new_n670), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(G1986), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT22), .B(G1981), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G29), .A2(G32), .ZN(new_n682));
  INV_X1    g257(.A(G129), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n632), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT92), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  AOI211_X1 g263(.A(new_n684), .B(new_n688), .C1(G105), .C2(new_n491), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n477), .A2(G141), .A3(new_n479), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT90), .Z(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n682), .B1(new_n692), .B2(G29), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT27), .B(G1996), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n491), .A2(G103), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  INV_X1    g275(.A(G139), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n699), .B1(new_n459), .B2(new_n700), .C1(new_n480), .C2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT89), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G29), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G29), .B2(G33), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(KEYINPUT23), .A3(G20), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n710));
  INV_X1    g285(.A(G20), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n712), .C1(new_n571), .C2(new_n708), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1956), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n696), .A2(new_n707), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n708), .A2(G19), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n549), .B2(new_n708), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1341), .Z(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2078), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n719), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT96), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT29), .ZN(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n705), .A2(new_n706), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n715), .A2(new_n718), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n693), .A2(new_n694), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(KEYINPUT24), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n719), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n719), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G2084), .Z(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G28), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G28), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(new_n741), .A3(new_n719), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n731), .A2(new_n732), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n726), .A2(new_n727), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n719), .A2(G26), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT87), .Z(new_n748));
  INV_X1    g323(.A(G128), .ZN(new_n749));
  INV_X1    g324(.A(G140), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n748), .B1(new_n749), .B2(new_n632), .C1(new_n480), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(G29), .ZN(new_n752));
  MUX2_X1   g327(.A(new_n745), .B(new_n752), .S(KEYINPUT28), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n755));
  NOR2_X1   g330(.A1(G286), .A2(new_n708), .ZN(new_n756));
  MUX2_X1   g331(.A(new_n755), .B(KEYINPUT94), .S(new_n756), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1966), .ZN(new_n758));
  NAND2_X1  g333(.A1(G171), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G5), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n754), .B(new_n758), .C1(G1961), .C2(new_n761), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n730), .A2(new_n743), .A3(new_n744), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n719), .A2(G25), .ZN(new_n764));
  OR2_X1    g339(.A1(G95), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n766));
  INV_X1    g341(.A(G119), .ZN(new_n767));
  INV_X1    g342(.A(G131), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n766), .B1(new_n767), .B2(new_n632), .C1(new_n480), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT81), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n719), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT83), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT35), .B(G1991), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT82), .Z(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n773), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G23), .ZN(new_n778));
  XNOR2_X1  g353(.A(G288), .B(KEYINPUT85), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n708), .A2(G6), .ZN(new_n783));
  INV_X1    g358(.A(G305), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n708), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT32), .B(G1981), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n782), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n794));
  MUX2_X1   g369(.A(G24), .B(G290), .S(G16), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT84), .B(G1986), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n793), .A2(KEYINPUT86), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n777), .A2(new_n798), .A3(KEYINPUT36), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT36), .B1(new_n777), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n708), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n612), .B2(new_n708), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n634), .A2(new_n719), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT95), .Z(new_n807));
  NAND4_X1  g382(.A1(new_n763), .A2(new_n801), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n761), .A2(G1961), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(G311));
  NAND2_X1  g386(.A1(G311), .A2(KEYINPUT97), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n808), .B2(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(G150));
  AOI22_X1  g390(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n497), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G55), .B2(new_n504), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n511), .A2(G93), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT99), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n612), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT39), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n548), .A2(new_n819), .A3(new_n818), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n820), .A2(new_n546), .A3(new_n547), .A4(new_n544), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n823), .B1(new_n831), .B2(G860), .ZN(G145));
  NAND2_X1  g407(.A1(new_n493), .A2(KEYINPUT100), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n489), .A2(G2105), .B1(G102), .B2(new_n491), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n486), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n692), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n751), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n751), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n703), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n703), .B(KEYINPUT101), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n839), .A2(new_n845), .A3(new_n840), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(G106), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n849));
  INV_X1    g424(.A(G130), .ZN(new_n850));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n849), .B1(new_n850), .B2(new_n632), .C1(new_n480), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n626), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n844), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n634), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n482), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n770), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  INV_X1    g437(.A(new_n860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n854), .A2(new_n856), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g441(.A(new_n621), .B(new_n830), .Z(new_n867));
  OAI211_X1 g442(.A(new_n571), .B(new_n600), .C1(new_n606), .C2(new_n610), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n604), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n571), .B1(new_n872), .B2(new_n600), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT41), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n611), .A2(G299), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n868), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT102), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n869), .A2(new_n873), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n867), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n867), .B2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n506), .B2(new_n515), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n499), .A2(KEYINPUT6), .A3(G651), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT6), .B1(new_n499), .B2(G651), .ZN(new_n888));
  OAI211_X1 g463(.A(G50), .B(G543), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT68), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n504), .A2(new_n495), .A3(G50), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n520), .B(G88), .C1(new_n887), .C2(new_n888), .ZN(new_n893));
  INV_X1    g468(.A(new_n513), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n520), .B2(G62), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n895), .B2(new_n497), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n892), .A2(KEYINPUT103), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G290), .B1(new_n886), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n892), .B2(new_n896), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n515), .A2(new_n885), .A3(new_n890), .A4(new_n891), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n589), .A4(new_n594), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n898), .A2(G305), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G305), .B1(new_n898), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n779), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND4_X1   g479(.A1(new_n589), .A2(new_n899), .A3(new_n900), .A4(new_n594), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n899), .A2(new_n900), .B1(new_n589), .B2(new_n594), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n784), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n779), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n898), .A2(G305), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI211_X1 g485(.A(KEYINPUT105), .B(KEYINPUT42), .C1(new_n904), .C2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n904), .A2(KEYINPUT104), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n904), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(KEYINPUT105), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n884), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n884), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n820), .A2(new_n596), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND2_X1  g501(.A1(G301), .A2(G168), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n530), .B(G286), .C1(new_n536), .C2(new_n537), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n830), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n828), .A2(new_n927), .A3(new_n829), .A4(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n878), .B2(new_n881), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n904), .A2(new_n910), .A3(KEYINPUT104), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n902), .A2(new_n903), .A3(new_n779), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n916), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n930), .A2(new_n931), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n880), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n934), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n939), .A4(new_n933), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n913), .B2(new_n914), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n937), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n933), .A2(new_n939), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(new_n939), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n938), .B1(new_n877), .B2(new_n874), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n944), .A2(new_n956), .A3(new_n957), .A4(new_n862), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n951), .A2(new_n957), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n944), .A2(new_n956), .A3(KEYINPUT43), .A4(new_n862), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n926), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT109), .B(new_n966), .C1(new_n961), .C2(new_n962), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(G397));
  NOR2_X1   g545(.A1(new_n837), .A2(G1384), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(G40), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(G290), .B(G1986), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n975), .A2(G1996), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n979), .B(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n751), .B(G2067), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n981), .A2(new_n692), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n692), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n976), .A2(G1996), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT111), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n770), .A2(new_n775), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n771), .A2(new_n776), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n976), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n971), .A2(new_n974), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT112), .B(G8), .Z(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(G305), .B(G1981), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT113), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n994), .B1(G1976), .B2(new_n779), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n837), .A2(new_n1007), .A3(G1384), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n486), .B2(new_n493), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n973), .B1(new_n1011), .B2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n790), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n833), .A2(new_n836), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n484), .B(KEYINPUT4), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1010), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n974), .B(new_n1015), .C1(new_n1019), .C2(KEYINPUT50), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(G2090), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1006), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT55), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n1017), .B2(new_n834), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n973), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n971), .B2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1014), .B1(G2090), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n993), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1024), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G288), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1002), .B(new_n1003), .C1(G1976), .C2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1005), .A2(new_n1025), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1019), .A2(new_n1007), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n974), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1039));
  INV_X1    g614(.A(G1966), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1020), .A2(G2084), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(new_n993), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G286), .A2(new_n993), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT121), .Z(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1044), .A2(KEYINPUT51), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1006), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1046), .B(KEYINPUT122), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1051), .A2(new_n1052), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1048), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT125), .B(G1961), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1020), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1012), .B(new_n1058), .C1(new_n1019), .C2(new_n1007), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(KEYINPUT126), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT126), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(G2078), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1039), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1068), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1037), .B1(new_n1055), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(G171), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n571), .B(KEYINPUT57), .ZN(new_n1073));
  INV_X1    g648(.A(G1956), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1029), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1009), .A2(new_n1012), .A3(new_n1076), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT61), .B(new_n1073), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n1079));
  INV_X1    g654(.A(G2067), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n971), .A2(new_n1079), .A3(new_n1080), .A4(new_n974), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1018), .A2(new_n974), .A3(new_n1010), .A4(new_n1080), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1020), .A2(new_n804), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(new_n1085), .A3(new_n1084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1078), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1093));
  NAND2_X1  g668(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(new_n1073), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1093), .B2(new_n1073), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n971), .B2(new_n974), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1098), .B(new_n1102), .C1(new_n1013), .C2(G1996), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n974), .B1(new_n1026), .B2(KEYINPUT45), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1008), .A2(new_n1104), .A3(G1996), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT118), .B1(new_n1105), .B2(new_n1101), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n549), .ZN(new_n1108));
  NAND2_X1  g683(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1107), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n549), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1092), .A2(new_n1097), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1093), .A2(new_n1073), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1093), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1073), .B(KEYINPUT117), .Z(new_n1115));
  AOI22_X1  g690(.A1(new_n1113), .A2(new_n612), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1009), .A2(new_n974), .A3(new_n1038), .A4(new_n1064), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1057), .B(new_n1117), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1118), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT127), .B1(new_n1118), .B2(G171), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1067), .B2(G301), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1112), .A2(new_n1116), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1071), .B1(G171), .B2(new_n1118), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1072), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1070), .B1(new_n1128), .B2(new_n1055), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1005), .A2(new_n1035), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1032), .A2(KEYINPUT115), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1022), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1044), .A2(G168), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1022), .A2(new_n1132), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1130), .A2(new_n1133), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT114), .B(KEYINPUT63), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1036), .B2(new_n1134), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1130), .A2(new_n1024), .A3(new_n1022), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1001), .A2(G1976), .A3(G288), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G305), .A2(G1981), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n995), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n978), .B(new_n991), .C1(new_n1129), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n987), .A2(new_n988), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n751), .A2(G2067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n975), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n981), .B(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n976), .B1(new_n984), .B2(new_n982), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT47), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n975), .A2(G1986), .A3(G290), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT48), .Z(new_n1157));
  AOI211_X1 g732(.A(new_n1149), .B(new_n1155), .C1(new_n991), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1146), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G401), .A2(G227), .ZN(new_n1161));
  AND2_X1   g735(.A1(new_n865), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g736(.A1(new_n1162), .A2(G319), .A3(new_n680), .A4(new_n961), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


