//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n462), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  XOR2_X1   g043(.A(KEYINPUT3), .B(G2104), .Z(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT65), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n477), .B2(G2105), .ZN(G160));
  NAND2_X1  g053(.A1(new_n465), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT66), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n472), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(new_n485), .B2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  INV_X1    g064(.A(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n484), .A2(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n465), .A2(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n465), .A2(new_n496), .A3(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT67), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT68), .B(G88), .Z(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(new_n499), .B1(G50), .B2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n504), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n503), .B2(new_n504), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT67), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT67), .A2(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT6), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n508), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(KEYINPUT69), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n516), .A2(G51), .A3(G543), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  OAI211_X1 g104(.A(G63), .B(G651), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n519), .B2(new_n520), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT70), .B(G89), .Z(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(G168));
  NAND4_X1  g112(.A1(new_n516), .A2(G52), .A3(G543), .A4(new_n521), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n532), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n541), .A2(new_n543), .B1(new_n509), .B2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n519), .A2(new_n520), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n513), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(G43), .A3(new_n521), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n532), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n533), .A2(G81), .B1(new_n554), .B2(new_n509), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n533), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n532), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n516), .A2(G53), .A3(G543), .A4(new_n521), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n550), .A2(new_n571), .A3(G53), .A4(new_n521), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n546), .A2(new_n509), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n542), .B1(new_n538), .B2(new_n539), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(G301));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n522), .A2(new_n535), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(new_n522), .B2(new_n535), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND4_X1  g158(.A1(new_n516), .A2(G49), .A3(G543), .A4(new_n521), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n502), .B1(new_n532), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n533), .B2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n532), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(new_n509), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n499), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n510), .B2(new_n593), .ZN(G305));
  NAND3_X1  g169(.A1(new_n550), .A2(G47), .A3(new_n521), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT73), .B(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n532), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n533), .A2(new_n596), .B1(new_n599), .B2(new_n509), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(G290));
  NAND4_X1  g176(.A1(new_n516), .A2(G54), .A3(G543), .A4(new_n521), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n502), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT10), .B1(new_n533), .B2(G92), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n602), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G284));
  OAI21_X1  g185(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G321));
  NOR2_X1   g186(.A1(G286), .A2(new_n608), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n573), .B(KEYINPUT74), .Z(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n608), .ZN(G297));
  AOI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n608), .ZN(G280));
  INV_X1    g190(.A(new_n607), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n556), .A2(new_n608), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n607), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n472), .A2(new_n466), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT13), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n465), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n490), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n484), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT75), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n635), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n652), .A3(new_n648), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(KEYINPUT77), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(KEYINPUT77), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT78), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n658), .B(new_n651), .C1(new_n654), .C2(new_n655), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT80), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n664), .A2(new_n666), .ZN(new_n672));
  INV_X1    g247(.A(new_n663), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n667), .B1(new_n673), .B2(new_n666), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n685), .B2(new_n691), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n694), .B(KEYINPUT81), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(KEYINPUT82), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n682), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(KEYINPUT82), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n696), .A2(new_n697), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n705), .A3(new_n681), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n701), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n701), .B2(new_n706), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n680), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n701), .A2(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(new_n702), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n701), .A2(new_n703), .A3(new_n706), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n711), .A2(new_n679), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(G229));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G129), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT88), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n715), .A2(G35), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n487), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n726), .A2(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n536), .A2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G21), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT90), .B(G1966), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n557), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G16), .B2(G19), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n733), .B(new_n739), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n735), .A2(G4), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n616), .B2(new_n735), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1348), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n740), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n747), .B1(new_n731), .B2(new_n732), .C1(new_n726), .C2(new_n727), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n743), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n715), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n485), .A2(G128), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n465), .A2(G140), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n490), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n715), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT85), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G33), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT86), .Z(new_n763));
  AND2_X1   g338(.A1(new_n472), .A2(G127), .ZN(new_n764));
  AND2_X1   g339(.A1(G115), .A2(G2104), .ZN(new_n765));
  OAI21_X1  g340(.A(G2105), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n490), .A2(G103), .A3(G2104), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(new_n465), .B2(G139), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n763), .B1(new_n772), .B2(new_n715), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT30), .B(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n777), .A2(new_n715), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n631), .B2(new_n715), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n775), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n715), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n715), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n782), .B(new_n786), .C1(new_n724), .C2(new_n725), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n737), .A2(new_n738), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n761), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT24), .ZN(new_n790));
  INV_X1    g365(.A(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G160), .B2(new_n715), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT87), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n735), .A2(G5), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G171), .B2(new_n735), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT91), .B(G1961), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n789), .B(new_n796), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT93), .B(KEYINPUT23), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n735), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n573), .B2(new_n735), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT94), .B(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n798), .B2(new_n800), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n749), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(G25), .A2(G29), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n465), .A2(G131), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n490), .ZN(new_n815));
  INV_X1    g390(.A(G119), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n484), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n817), .B2(new_n715), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT83), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G290), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G16), .B2(G24), .ZN(new_n824));
  INV_X1    g399(.A(G1986), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n584), .A2(new_n587), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n735), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n735), .B2(G23), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT33), .B(G1976), .Z(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n735), .A2(G22), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G166), .B2(new_n735), .ZN(new_n837));
  INV_X1    g412(.A(G1971), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G6), .A2(G16), .ZN(new_n840));
  INV_X1    g415(.A(new_n592), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n593), .A2(new_n510), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n840), .B1(new_n843), .B2(G16), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT32), .B(G1981), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n834), .A2(new_n835), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n828), .B1(new_n847), .B2(KEYINPUT34), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT84), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n811), .B1(new_n852), .B2(new_n854), .ZN(G311));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n810), .ZN(G150));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  INV_X1    g433(.A(G67), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n532), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n533), .A2(G93), .B1(new_n860), .B2(new_n509), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n516), .A2(G55), .A3(G543), .A4(new_n521), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  INV_X1    g440(.A(new_n863), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n557), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(KEYINPUT96), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n556), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n616), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G860), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(KEYINPUT98), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT98), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n865), .B1(new_n882), .B2(new_n883), .ZN(G145));
  NAND2_X1  g459(.A1(new_n495), .A2(new_n497), .ZN(new_n885));
  INV_X1    g460(.A(new_n493), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n756), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n485), .A2(G130), .B1(G142), .B2(new_n465), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(KEYINPUT101), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n892), .A2(new_n490), .A3(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n490), .B2(G118), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n893), .B(new_n894), .C1(KEYINPUT101), .C2(new_n890), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n889), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n888), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n817), .B(KEYINPUT102), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n624), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n772), .B(new_n721), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n487), .B(new_n631), .Z(new_n908));
  XNOR2_X1  g483(.A(G160), .B(KEYINPUT99), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n910), .B2(new_n907), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g488(.A1(new_n863), .A2(new_n608), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n872), .B(new_n620), .ZN(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(new_n607), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n616), .A2(new_n573), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n616), .A2(new_n573), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n616), .A2(new_n573), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT41), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n923), .A3(new_n917), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(KEYINPUT103), .A3(KEYINPUT41), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n915), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT104), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G303), .B(G290), .ZN(new_n930));
  XNOR2_X1  g505(.A(G288), .B(G305), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT42), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n919), .A2(KEYINPUT104), .A3(new_n928), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n934), .B(new_n935), .Z(new_n936));
  OAI21_X1  g511(.A(new_n914), .B1(new_n936), .B2(new_n608), .ZN(G295));
  OAI21_X1  g512(.A(new_n914), .B1(new_n936), .B2(new_n608), .ZN(G331));
  NAND3_X1  g513(.A1(G301), .A2(KEYINPUT105), .A3(G168), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n541), .A2(new_n543), .ZN(new_n940));
  NAND3_X1  g515(.A1(G286), .A2(new_n940), .A3(new_n575), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(G301), .B2(G168), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n872), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n868), .A2(new_n871), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G171), .B2(new_n536), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n945), .A2(new_n947), .A3(new_n941), .A4(new_n939), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n920), .A2(new_n921), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n944), .A2(new_n926), .A3(new_n948), .A4(new_n927), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n932), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n957), .A3(new_n923), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n918), .A2(new_n960), .A3(KEYINPUT41), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n956), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n948), .A3(new_n944), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n932), .B1(new_n963), .B2(new_n951), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n932), .B1(new_n951), .B2(new_n952), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(G37), .ZN(new_n970));
  INV_X1    g545(.A(new_n932), .ZN(new_n971));
  AND4_X1   g546(.A1(new_n927), .A2(new_n944), .A3(new_n926), .A4(new_n948), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n918), .B1(new_n944), .B2(new_n948), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT106), .A3(new_n954), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(new_n975), .A3(new_n976), .A4(new_n953), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n955), .C2(new_n964), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n967), .A2(new_n977), .A3(KEYINPUT44), .A4(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n955), .A2(new_n964), .A3(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(new_n975), .A3(new_n953), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT43), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(KEYINPUT44), .B2(new_n982), .ZN(G397));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n887), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT111), .B1(new_n887), .B2(new_n984), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n987), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n471), .A2(new_n474), .B1(G113), .B2(G2104), .ZN(new_n990));
  OAI211_X1 g565(.A(G40), .B(new_n467), .C1(new_n990), .C2(new_n490), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n756), .B(new_n760), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n996), .B2(new_n722), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(G1996), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n994), .A2(new_n997), .B1(new_n722), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n820), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n817), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n817), .A2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n993), .ZN(new_n1005));
  XNOR2_X1  g580(.A(G290), .B(G1986), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT124), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n536), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT125), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1008), .B(KEYINPUT51), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n992), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n738), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n887), .A2(new_n1019), .A3(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n992), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(G2084), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n1011), .C1(new_n1022), .C2(new_n536), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1009), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1022), .A2(new_n1024), .B1(new_n1008), .B2(KEYINPUT51), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1010), .A2(KEYINPUT51), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n992), .A2(new_n1020), .A3(new_n1018), .ZN(new_n1027));
  INV_X1    g602(.A(G2084), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1027), .A2(new_n1028), .B1(new_n1016), .B2(new_n738), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1009), .B(new_n1026), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1023), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G166), .A2(new_n1030), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1037), .B2(KEYINPUT55), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n992), .A2(new_n1013), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1027), .A2(new_n732), .B1(new_n1041), .B2(new_n838), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1042), .B2(new_n1030), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n829), .A2(G1976), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n887), .A2(new_n1014), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1044), .B(G8), .C1(new_n991), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  NAND4_X1  g622(.A1(G160), .A2(G40), .A3(new_n1014), .A4(new_n887), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(G8), .A3(new_n1044), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  INV_X1    g627(.A(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(new_n842), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n592), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n843), .A2(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1048), .A2(new_n1057), .A3(new_n1060), .A4(G8), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1047), .A2(new_n1051), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1043), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1021), .B2(G2090), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1041), .A2(new_n838), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n991), .B1(new_n1045), .B2(KEYINPUT50), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT113), .A3(new_n732), .A4(new_n1020), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1039), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(G171), .B(KEYINPUT54), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n992), .A2(new_n1013), .A3(new_n1040), .A4(new_n785), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n1075), .B1(new_n1021), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n490), .B1(new_n477), .B2(KEYINPUT126), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(KEYINPUT126), .B2(new_n477), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1074), .A2(G2078), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n467), .A2(G40), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1040), .A3(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1073), .B(new_n1077), .C1(new_n989), .C2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n992), .A2(new_n1013), .A3(new_n1015), .A4(new_n1080), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1085), .B2(new_n1073), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1072), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n992), .A2(new_n1013), .A3(new_n1040), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(G2072), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1088), .A2(new_n1090), .B1(new_n1021), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n568), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n1093), .B2(KEYINPUT119), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(new_n573), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1045), .A2(new_n991), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1021), .A2(new_n1098), .B1(new_n760), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n607), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n992), .A2(new_n1013), .A3(new_n1040), .A4(new_n1090), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1027), .B2(G1956), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT121), .B(new_n1102), .C1(new_n1027), .C2(G1956), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1095), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1105), .A2(KEYINPUT122), .A3(new_n1107), .A4(new_n1106), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1097), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT123), .B(G1996), .Z(new_n1113));
  NAND4_X1  g688(.A1(new_n992), .A2(new_n1013), .A3(new_n1040), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1045), .B2(new_n991), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n557), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n557), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1119), .A2(new_n1121), .B1(new_n1100), .B2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1100), .A2(new_n607), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1101), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1096), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1092), .A2(new_n1126), .A3(new_n1095), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n1123), .A2(new_n1125), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1087), .B1(new_n1112), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1132));
  AOI21_X1  g707(.A(G301), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1071), .A3(new_n1063), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1033), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1029), .A2(new_n1030), .A3(G286), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1071), .A4(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1071), .A2(new_n1136), .A3(new_n1043), .A4(new_n1062), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1071), .A2(new_n1136), .A3(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1069), .A2(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1039), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT118), .B1(new_n1145), .B2(new_n1062), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1047), .A2(new_n1061), .A3(new_n1051), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1147), .B(new_n1148), .C1(new_n1144), .C2(new_n1039), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1143), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1142), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1071), .A2(new_n1043), .A3(new_n1062), .A4(new_n1133), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(KEYINPUT62), .B2(new_n1032), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1062), .A2(new_n1069), .A3(G8), .A4(new_n1070), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1099), .A2(new_n1030), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1061), .A2(new_n1049), .A3(new_n829), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1056), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT115), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1154), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1153), .A2(KEYINPUT62), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1151), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1007), .B1(new_n1135), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n998), .B(KEYINPUT46), .Z(new_n1165));
  INV_X1    g740(.A(new_n995), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n994), .B1(new_n721), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n993), .A2(G1986), .A3(G290), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1170), .A2(new_n1171), .B1(new_n1004), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n999), .A2(new_n1001), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(G2067), .B2(new_n756), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(new_n994), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1164), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g753(.A1(G227), .A2(new_n459), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n657), .B2(new_n659), .ZN(new_n1181));
  NAND4_X1  g755(.A1(new_n1181), .A2(new_n709), .A3(new_n713), .A4(new_n912), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n982), .A2(new_n1182), .ZN(G308));
  OR2_X1    g757(.A1(new_n982), .A2(new_n1182), .ZN(G225));
endmodule


