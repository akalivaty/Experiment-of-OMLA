//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(new_n448), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(new_n469), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n464), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n488), .B1(new_n487), .B2(new_n486), .C1(G112), .C2(new_n469), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n467), .A2(new_n482), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT71), .B1(new_n475), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n467), .A2(new_n494), .A3(new_n478), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(G136), .B2(new_n496), .ZN(G162));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n473), .B2(new_n474), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G138), .B1(new_n473), .B2(new_n474), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n504), .B2(new_n482), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n467), .A2(new_n469), .A3(new_n506), .A4(G138), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n516), .A2(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n512), .B1(new_n526), .B2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n516), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n519), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n511), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n516), .A2(new_n541), .B1(new_n522), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n540), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n516), .A2(new_n546), .B1(new_n522), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n509), .A2(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n511), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n548), .B1(new_n552), .B2(KEYINPUT74), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n522), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n515), .A2(new_n509), .A3(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(G91), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n565), .A2(KEYINPUT80), .A3(G91), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT81), .B(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n534), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n513), .B2(new_n514), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(G53), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n576), .A2(KEYINPUT78), .A3(G53), .A4(new_n577), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT9), .B1(new_n516), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n574), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND3_X1  g161(.A1(new_n565), .A2(G87), .A3(new_n566), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n576), .B2(G49), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n534), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G48), .B2(new_n576), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n565), .A2(G86), .A3(new_n566), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n576), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI221_X1 g175(.A(new_n598), .B1(new_n599), .B2(new_n522), .C1(new_n600), .C2(new_n511), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n576), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(G54), .B1(new_n576), .B2(KEYINPUT82), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n604), .A2(new_n605), .B1(new_n511), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n565), .A2(new_n566), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n608), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n607), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n602), .B1(new_n613), .B2(G868), .ZN(G284));
  XOR2_X1   g189(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g200(.A(new_n491), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n496), .A2(G135), .B1(G123), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n469), .A2(new_n628), .A3(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n469), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n627), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n467), .A2(new_n470), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT13), .B(G2100), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n647), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(new_n655), .A3(G14), .ZN(G401));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT87), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT89), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n662), .A3(new_n660), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n658), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n662), .B1(new_n670), .B2(new_n661), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  XNOR2_X1  g267(.A(KEYINPUT90), .B(G29), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  OAI221_X1 g270(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n496), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n626), .A2(G119), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT92), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n695), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT93), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT33), .B(G1976), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  MUX2_X1   g289(.A(G6), .B(G305), .S(G16), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XOR2_X1   g291(.A(new_n715), .B(new_n716), .Z(new_n717));
  NOR3_X1   g292(.A1(new_n708), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  MUX2_X1   g296(.A(G24), .B(G290), .S(G16), .Z(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1986), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n705), .A2(new_n724), .A3(KEYINPUT36), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT36), .B1(new_n705), .B2(new_n724), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT24), .B(G34), .ZN(new_n728));
  AOI22_X1  g303(.A1(G160), .A2(G29), .B1(new_n693), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G2084), .ZN(new_n730));
  NOR2_X1   g305(.A1(G171), .A2(new_n709), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G5), .B2(new_n709), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  OAI22_X1  g308(.A1(new_n732), .A2(new_n733), .B1(new_n632), .B2(new_n693), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n730), .B(new_n734), .C1(new_n733), .C2(new_n732), .ZN(new_n735));
  NOR2_X1   g310(.A1(G168), .A2(new_n709), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n709), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT96), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G28), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n745), .B1(new_n743), .B2(G28), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n729), .B2(G2084), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n742), .A2(G33), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n496), .A2(G139), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n755), .C1(new_n469), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n749), .B1(new_n750), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n737), .A2(new_n738), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n735), .A2(new_n740), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n742), .A2(G32), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT26), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(G105), .B2(new_n470), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n491), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n496), .B2(G141), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n742), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G162), .A2(new_n694), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G35), .B2(new_n694), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT29), .ZN(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n774), .B1(new_n750), .B2(new_n758), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n693), .A2(G27), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT99), .Z(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n693), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT100), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  INV_X1    g359(.A(new_n777), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G2090), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n762), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n693), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n496), .A2(G140), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n469), .A2(G116), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n626), .A2(G128), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(new_n742), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n709), .A2(G19), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n557), .B2(new_n709), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1341), .ZN(new_n803));
  NOR2_X1   g378(.A1(G4), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n613), .B2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n803), .B1(new_n805), .B2(G1348), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n800), .B(new_n806), .C1(G1348), .C2(new_n805), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n709), .A2(G20), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT23), .Z(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n787), .A2(new_n808), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n727), .A2(new_n814), .ZN(G311));
  INV_X1    g390(.A(G311), .ZN(G150));
  AOI22_X1  g391(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n511), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n516), .A2(new_n819), .B1(new_n522), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n613), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n557), .A2(KEYINPUT102), .A3(new_n822), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n822), .A2(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n822), .A2(KEYINPUT102), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n556), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n828), .B(new_n833), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n823), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n825), .B1(new_n836), .B2(new_n837), .ZN(G145));
  NAND2_X1  g413(.A1(new_n505), .A2(new_n507), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n500), .B1(new_n465), .B2(new_n466), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n478), .A2(G114), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n499), .A2(KEYINPUT104), .A3(new_n502), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT103), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n841), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n796), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n637), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n496), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n626), .A2(G130), .ZN(new_n856));
  OAI221_X1 g431(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n701), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n701), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n757), .B(new_n771), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n861), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n854), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n853), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n632), .B(G160), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n867), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n879));
  XNOR2_X1  g454(.A(G288), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G305), .ZN(new_n881));
  XOR2_X1   g456(.A(G303), .B(G290), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n833), .B(new_n622), .Z(new_n886));
  INV_X1    g461(.A(new_n613), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n617), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n613), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT105), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n888), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n888), .B2(new_n889), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n886), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n833), .B(new_n622), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n890), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n885), .B1(new_n901), .B2(KEYINPUT108), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(KEYINPUT108), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n885), .A3(KEYINPUT108), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G868), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n822), .A2(G868), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(G295));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n911), .A3(new_n909), .ZN(new_n912));
  INV_X1    g487(.A(G868), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n904), .B2(new_n905), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT109), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(G331));
  OAI21_X1  g491(.A(G168), .B1(G301), .B2(KEYINPUT110), .ZN(new_n917));
  NAND2_X1  g492(.A1(G301), .A2(KEYINPUT110), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n917), .B(new_n918), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n833), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(new_n891), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n896), .B2(new_n920), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(new_n883), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n922), .B2(new_n883), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n896), .A2(new_n920), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n883), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n876), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n890), .A2(new_n893), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n920), .B(new_n931), .C1(KEYINPUT41), .C2(new_n890), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n883), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n925), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n930), .B1(new_n923), .B2(new_n924), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n929), .A2(KEYINPUT43), .A3(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n938), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n849), .A2(new_n850), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT103), .B1(new_n505), .B2(new_n507), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n471), .A2(G40), .A3(new_n483), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n796), .B(new_n799), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT111), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(new_n771), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(G1996), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n954), .A3(new_n771), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n701), .A2(new_n704), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n701), .A2(new_n704), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n947), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT48), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n955), .A3(new_n959), .A4(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n951), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n947), .A2(new_n954), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n964), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n956), .B(KEYINPUT127), .Z(new_n972));
  NAND3_X1  g547(.A1(new_n953), .A2(new_n955), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n797), .A2(new_n799), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n948), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1956), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n851), .B2(new_n940), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n471), .A2(G40), .A3(new_n483), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n505), .A2(new_n507), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n940), .B1(new_n981), .B2(new_n503), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n977), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n946), .B1(new_n982), .B2(new_n944), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT45), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT56), .B(G2072), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n569), .A2(new_n570), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n573), .A2(G651), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(KEYINPUT57), .A3(new_n584), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT120), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n574), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n584), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n580), .A2(new_n583), .A3(new_n997), .A4(new_n581), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n584), .A2(KEYINPUT119), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n574), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n994), .A2(new_n995), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n989), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n995), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n996), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1004), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n978), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n851), .A2(KEYINPUT112), .A3(new_n978), .A4(new_n940), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G164), .A2(G1384), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT113), .B1(new_n1013), .B2(new_n978), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n982), .A2(new_n1015), .A3(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n946), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1348), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n851), .A2(new_n980), .A3(new_n940), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2067), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n989), .A2(new_n1001), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n887), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1007), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(KEYINPUT60), .A3(new_n1023), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT60), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1348), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n1022), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n613), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n989), .A2(new_n1001), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n1025), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1020), .A2(KEYINPUT60), .A3(new_n887), .A4(new_n1023), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n985), .A2(new_n954), .A3(new_n986), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n985), .A2(KEYINPUT122), .A3(new_n986), .A4(new_n954), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT58), .B(G1341), .Z(new_n1042));
  NAND2_X1  g617(.A1(new_n1021), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n557), .ZN(new_n1045));
  NAND2_X1  g620(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1044), .A2(KEYINPUT123), .A3(KEYINPUT59), .A4(new_n557), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT61), .B1(new_n989), .B2(new_n1001), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1047), .B(new_n1048), .C1(new_n1007), .C2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1027), .B1(new_n1037), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1012), .A2(new_n1017), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n1054));
  NOR3_X1   g629(.A1(G164), .A2(new_n944), .A3(G1384), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT118), .B(G1966), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n849), .A2(new_n850), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1384), .B1(new_n1059), .B2(new_n841), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n980), .B(new_n1056), .C1(new_n1060), .C2(KEYINPUT45), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1061), .B2(new_n738), .ZN(new_n1062));
  OAI211_X1 g637(.A(G168), .B(new_n1053), .C1(new_n1057), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1053), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(G286), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1054), .A2(new_n986), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2078), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n986), .A2(new_n1074), .A3(new_n980), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1071), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1961), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1070), .B1(new_n1080), .B2(G301), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1079), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n946), .B(new_n1055), .C1(new_n943), .C2(new_n944), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1083), .A2(new_n1072), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(new_n1070), .A3(G301), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n587), .A2(G1976), .A3(new_n590), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(new_n1021), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  INV_X1    g669(.A(G1976), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(G288), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(G8), .A3(new_n1021), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n594), .A2(G651), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n576), .A2(G48), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n515), .A2(new_n509), .A3(G86), .ZN(new_n1101));
  OAI21_X1  g676(.A(G1981), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1103));
  INV_X1    g678(.A(G1981), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n595), .A2(new_n596), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1102), .A2(new_n1105), .A3(KEYINPUT115), .A4(KEYINPUT49), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(G8), .A3(new_n1021), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1094), .A2(new_n1097), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1094), .A2(KEYINPUT117), .A3(new_n1110), .A4(new_n1097), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n979), .A2(new_n983), .A3(G2090), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1971), .B1(new_n985), .B2(new_n986), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n946), .B1(new_n1013), .B2(new_n978), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n778), .B(new_n1120), .C1(new_n1060), .C2(new_n978), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n985), .A2(new_n986), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1121), .B(KEYINPUT116), .C1(new_n1122), .C2(G1971), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G303), .A2(G8), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT55), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1018), .A2(G2090), .B1(G1971), .B2(new_n1122), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1126), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(G8), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1082), .A2(G301), .A3(new_n1084), .ZN(new_n1132));
  OAI21_X1  g707(.A(G171), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT54), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1051), .A2(new_n1069), .A3(new_n1090), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1068), .A2(new_n1064), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1066), .B1(new_n1063), .B2(G8), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1065), .B(new_n1140), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1131), .A2(new_n1086), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1110), .A2(new_n1095), .A3(new_n711), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1105), .ZN(new_n1145));
  OAI211_X1 g720(.A(G8), .B(new_n1021), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1130), .B2(new_n1111), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  AND2_X1   g723(.A1(G168), .A2(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1067), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1131), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1128), .A2(G8), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1126), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1111), .A2(new_n1148), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1147), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1136), .A2(new_n1143), .A3(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n947), .B1(new_n960), .B2(new_n1159), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1160), .A2(new_n953), .A3(new_n955), .A4(new_n959), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1158), .A2(KEYINPUT126), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT126), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n976), .B1(new_n1162), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(new_n461), .ZN(new_n1166));
  NOR4_X1   g740(.A1(G229), .A2(new_n1166), .A3(G401), .A4(G227), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n877), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g742(.A1(new_n938), .A2(new_n1168), .ZN(G308));
  INV_X1    g743(.A(G308), .ZN(G225));
endmodule


