//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT77), .Z(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT66), .ZN(new_n195));
  OAI21_X1  g009(.A(G143), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G143), .Z(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G146), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n200), .A2(new_n194), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n194), .A2(KEYINPUT66), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n192), .A2(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT65), .A2(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT65), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(G146), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G128), .A3(new_n197), .ZN(new_n212));
  OAI21_X1  g026(.A(G128), .B1(new_n207), .B2(new_n197), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT71), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n194), .A3(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n205), .A2(new_n206), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n224), .B1(new_n221), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT78), .B1(new_n223), .B2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n223), .A2(KEYINPUT78), .A3(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n191), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n211), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n210), .A2(G146), .ZN(new_n238));
  AND4_X1   g052(.A1(G128), .A2(new_n238), .A3(new_n196), .A4(new_n197), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n234), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT10), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT67), .A2(G134), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n243), .A2(new_n246), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT68), .A2(G131), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(G137), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n247), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n250), .B(new_n251), .C1(new_n254), .C2(new_n243), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n243), .B1(new_n252), .B2(new_n253), .ZN(new_n256));
  OAI211_X1 g070(.A(KEYINPUT68), .B(G131), .C1(new_n256), .C2(new_n249), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OR3_X1    g073(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n217), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n238), .A2(new_n196), .A3(new_n259), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n225), .A2(new_n226), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n235), .A2(new_n242), .A3(new_n258), .A4(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n204), .A2(new_n212), .A3(new_n218), .A4(new_n233), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n240), .ZN(new_n273));
  INV_X1    g087(.A(new_n258), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT12), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n276));
  AOI211_X1 g090(.A(new_n276), .B(new_n258), .C1(new_n272), .C2(new_n240), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n271), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g093(.A(G227), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n279), .B(new_n281), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n235), .A2(new_n242), .A3(new_n270), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n274), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n271), .A3(new_n282), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(G469), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(G469), .A2(G902), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT79), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n274), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n276), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n273), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT80), .B1(new_n275), .B2(new_n277), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n271), .A2(new_n282), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT81), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n286), .A2(new_n271), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n283), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n190), .B1(new_n292), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n219), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n265), .A2(new_n312), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G224), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT7), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n313), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(G110), .B(G122), .Z(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT72), .B(G116), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT2), .B(G113), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n323), .A3(G116), .ZN(new_n330));
  OAI211_X1 g144(.A(G113), .B(new_n330), .C1(new_n326), .C2(new_n329), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n234), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n234), .B1(new_n328), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n322), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n319), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n326), .B(new_n327), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n269), .A2(new_n337), .A3(new_n267), .ZN(new_n338));
  INV_X1    g152(.A(new_n320), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n314), .B1(new_n219), .B2(new_n312), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n318), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n308), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT84), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n332), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n320), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n317), .B(KEYINPUT82), .Z(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n341), .A2(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n351), .A3(new_n320), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n308), .C1(new_n336), .C2(new_n342), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT85), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n344), .A2(new_n360), .A3(new_n353), .A4(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT86), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n364));
  OAI21_X1  g178(.A(G214), .B1(G237), .B2(G902), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n365), .A3(new_n363), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT87), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n311), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G131), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n256), .B2(new_n249), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n246), .A2(new_n248), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G137), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n247), .A2(G134), .ZN(new_n374));
  OAI21_X1  g188(.A(G131), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n219), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n266), .A2(new_n257), .A3(new_n255), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n258), .A2(new_n265), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n371), .A2(new_n381), .A3(new_n375), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n371), .B2(new_n375), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n384), .B2(new_n219), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n337), .B(new_n379), .C1(new_n385), .C2(KEYINPUT30), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n316), .A3(G210), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT27), .Z(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT26), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n226), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n380), .B1(new_n219), .B2(new_n376), .ZN(new_n392));
  INV_X1    g206(.A(new_n337), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n386), .A2(KEYINPUT73), .A3(new_n391), .A4(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(KEYINPUT31), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT31), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n394), .B(KEYINPUT28), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n385), .A2(new_n393), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n391), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G472), .A2(G902), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT32), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT32), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n399), .B2(new_n401), .ZN(new_n411));
  INV_X1    g225(.A(new_n408), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n377), .A2(new_n378), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n337), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n394), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT28), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT74), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n414), .A2(new_n337), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n419), .A2(KEYINPUT28), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n421), .A3(KEYINPUT28), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n424));
  INV_X1    g238(.A(new_n391), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(KEYINPUT28), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n420), .A2(new_n391), .A3(new_n404), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n424), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n386), .A2(new_n394), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n391), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n308), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G472), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n409), .A2(new_n413), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(new_n308), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT23), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n323), .B2(G128), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n438), .B(new_n439), .C1(G119), .C2(new_n191), .ZN(new_n440));
  XNOR2_X1  g254(.A(G119), .B(G128), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT24), .B(G110), .Z(new_n442));
  OAI22_X1  g256(.A1(new_n440), .A2(G110), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT16), .ZN(new_n445));
  OR3_X1    g259(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(G146), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n216), .A2(new_n444), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n440), .A2(G110), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT75), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n442), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n445), .A2(G146), .A3(new_n446), .ZN(new_n455));
  AOI21_X1  g269(.A(G146), .B1(new_n445), .B2(new_n446), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT22), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G137), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n458), .B(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n463), .A2(G902), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n458), .B(new_n461), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n308), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n436), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n436), .A2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G116), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(KEYINPUT72), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n325), .A2(KEYINPUT14), .A3(new_n477), .ZN(new_n484));
  OAI21_X1  g298(.A(G107), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n210), .A2(G128), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(G128), .B2(new_n202), .ZN(new_n488));
  INV_X1    g302(.A(new_n372), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n487), .B(new_n372), .C1(G128), .C2(new_n202), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT90), .B1(new_n481), .B2(new_n475), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n476), .C1(new_n325), .C2(new_n477), .ZN(new_n495));
  AOI21_X1  g309(.A(G107), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G107), .C1(new_n483), .C2(new_n484), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n486), .A2(new_n492), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n210), .A2(new_n501), .A3(G128), .ZN(new_n502));
  OAI211_X1 g316(.A(G134), .B(new_n502), .C1(new_n488), .C2(new_n501), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n493), .A2(new_n495), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n223), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n503), .B(new_n491), .C1(new_n505), .C2(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n187), .A2(G217), .A3(new_n316), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n308), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(KEYINPUT92), .A3(new_n308), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  MUX2_X1   g333(.A(new_n515), .B(new_n517), .S(new_n519), .Z(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(G952), .A3(new_n316), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G475), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n202), .A2(new_n387), .A3(new_n316), .A4(G214), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n387), .A2(new_n316), .A3(G214), .ZN(new_n529));
  OAI211_X1 g343(.A(G131), .B(new_n528), .C1(new_n210), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n528), .B1(new_n210), .B2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n370), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n530), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n457), .B(new_n532), .C1(KEYINPUT17), .C2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n221), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n533), .B1(new_n539), .B2(new_n370), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n448), .B1(new_n194), .B2(new_n444), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n540), .B(new_n541), .C1(new_n539), .C2(new_n530), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n538), .B1(new_n536), .B2(new_n542), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n527), .B1(new_n545), .B2(new_n308), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n444), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n312), .A2(G140), .ZN(new_n550));
  INV_X1    g364(.A(G140), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G125), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT19), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n553), .A3(new_n216), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n447), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n447), .A3(KEYINPUT88), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n535), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n538), .B1(new_n559), .B2(new_n542), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n527), .B(new_n308), .C1(new_n543), .C2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT89), .B1(new_n561), .B2(KEYINPUT20), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(KEYINPUT20), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n561), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n547), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n520), .A2(new_n526), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n369), .A2(new_n434), .A3(new_n473), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n407), .A2(new_n308), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n411), .B2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n292), .A2(new_n309), .ZN(new_n577));
  INV_X1    g391(.A(new_n190), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n473), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n570), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n190), .B(new_n472), .C1(new_n292), .C2(new_n309), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT94), .A3(new_n574), .A4(new_n575), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n365), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n359), .B2(new_n361), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n590));
  INV_X1    g404(.A(new_n511), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n510), .B1(new_n500), .B2(new_n506), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n509), .A2(new_n587), .A3(new_n588), .A4(new_n511), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(G478), .A3(new_n308), .ZN(new_n596));
  AOI21_X1  g410(.A(G478), .B1(new_n512), .B2(new_n308), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n566), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n586), .A2(new_n526), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  NAND3_X1  g418(.A1(new_n585), .A2(new_n520), .A3(new_n525), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n547), .A2(KEYINPUT96), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT20), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n558), .A2(new_n535), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT88), .B1(new_n554), .B2(new_n447), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n542), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n538), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(new_n613));
  AOI21_X1  g427(.A(G475), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n607), .B1(new_n614), .B2(new_n308), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n563), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n546), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n606), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n605), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n583), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT97), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT35), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n223), .ZN(G9));
  AOI21_X1  g438(.A(new_n573), .B1(new_n407), .B2(new_n308), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n411), .A2(G902), .A3(new_n572), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n462), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n458), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n470), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n469), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n369), .A2(new_n567), .A3(new_n627), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT37), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(G110), .Z(G12));
  INV_X1    g448(.A(new_n631), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n586), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n520), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n522), .B(KEYINPUT98), .Z(new_n638));
  OR2_X1    g452(.A1(new_n524), .A2(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n606), .A2(new_n616), .A3(new_n618), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n434), .A2(new_n310), .A3(new_n636), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  XOR2_X1   g458(.A(new_n640), .B(KEYINPUT39), .Z(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n310), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n520), .A2(new_n566), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n362), .A2(new_n363), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n362), .A2(KEYINPUT38), .A3(new_n363), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n648), .A2(new_n365), .A3(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n397), .A2(new_n398), .B1(new_n425), .B2(new_n416), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n656), .B2(G902), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n409), .A2(new_n413), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n635), .C1(KEYINPUT40), .C2(new_n647), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n210), .ZN(G45));
  NAND3_X1  g475(.A1(new_n566), .A2(new_n599), .A3(new_n640), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n434), .A2(new_n310), .A3(new_n664), .A4(new_n636), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT100), .B(G146), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G48));
  NAND2_X1  g481(.A1(new_n306), .A2(new_n308), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G469), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n578), .A3(new_n309), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n434), .A2(new_n671), .A3(new_n473), .A4(new_n601), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND4_X1  g488(.A1(new_n434), .A2(new_n671), .A3(new_n473), .A4(new_n620), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NAND4_X1  g490(.A1(new_n434), .A2(new_n671), .A3(new_n567), .A4(new_n636), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NAND3_X1  g492(.A1(new_n614), .A2(new_n607), .A3(new_n308), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n615), .B2(KEYINPUT89), .ZN(new_n680));
  INV_X1    g494(.A(new_n565), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n546), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n670), .A2(new_n605), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n423), .A2(new_n425), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n402), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n408), .B(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n411), .B2(G902), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n683), .A2(new_n684), .A3(new_n473), .A4(new_n690), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n585), .A2(new_n520), .A3(new_n525), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n692), .A2(new_n695), .A3(new_n566), .A4(new_n578), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n688), .A2(new_n689), .A3(new_n473), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT103), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n477), .ZN(G24));
  AND4_X1   g515(.A1(new_n578), .A2(new_n669), .A3(new_n309), .A4(new_n585), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n690), .A2(new_n631), .A3(new_n702), .A4(new_n664), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  AOI21_X1  g518(.A(KEYINPUT32), .B1(new_n407), .B2(new_n408), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n411), .A2(new_n410), .A3(new_n412), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT104), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n413), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n433), .A3(new_n709), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n283), .A2(new_n278), .B1(new_n299), .B2(new_n286), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(G902), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n190), .B1(new_n309), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n584), .B1(new_n362), .B2(new_n363), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n664), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n710), .A2(new_n715), .A3(new_n473), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n434), .A2(new_n473), .A3(new_n713), .A4(new_n714), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n664), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT105), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND2_X1  g537(.A1(new_n718), .A2(new_n642), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  AOI21_X1  g539(.A(KEYINPUT45), .B1(new_n284), .B2(new_n287), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n726), .B2(new_n307), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(G469), .C1(new_n711), .C2(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n289), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n693), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n289), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n190), .B(new_n645), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n597), .B1(new_n738), .B2(G478), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n566), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n682), .A2(new_n599), .A3(KEYINPUT43), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n631), .B(new_n742), .C1(new_n625), .C2(new_n626), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n635), .B1(new_n574), .B2(new_n575), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(KEYINPUT44), .A3(new_n742), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n736), .A2(new_n745), .A3(new_n714), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT107), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  AND3_X1   g564(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n289), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n731), .B2(new_n289), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n751), .A2(new_n752), .A3(new_n693), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT47), .B1(new_n753), .B2(new_n190), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n664), .A2(new_n714), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n434), .A2(new_n473), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n732), .A2(new_n733), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n309), .A3(new_n735), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n578), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT108), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n551), .ZN(G42));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n409), .A2(new_n413), .A3(new_n657), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n650), .A2(new_n365), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n670), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n472), .A2(new_n522), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n682), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n769), .B2(new_n599), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n695), .A2(new_n578), .A3(new_n714), .ZN(new_n771));
  INV_X1    g585(.A(new_n768), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n658), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n682), .A4(new_n739), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n638), .B1(new_n740), .B2(new_n741), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n671), .A2(new_n714), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n631), .A3(new_n690), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n695), .A2(KEYINPUT113), .A3(new_n584), .A4(new_n578), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n669), .A2(new_n584), .A3(new_n578), .A4(new_n309), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n473), .A2(new_n776), .A3(new_n689), .A4(new_n688), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n652), .A2(new_n653), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AND4_X1   g600(.A1(KEYINPUT50), .A2(new_n783), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n785), .B1(new_n779), .B2(new_n782), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT50), .B1(new_n788), .B2(new_n784), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n778), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n775), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n695), .A2(new_n190), .ZN(new_n792));
  INV_X1    g606(.A(new_n760), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n759), .B1(new_n758), .B2(new_n578), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n784), .A2(new_n714), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n791), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n778), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n788), .A2(new_n784), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n788), .A2(KEYINPUT50), .A3(new_n784), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n770), .A2(new_n774), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(KEYINPUT51), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n710), .A2(new_n473), .A3(new_n777), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(G952), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n813), .B(G953), .C1(new_n784), .C2(new_n702), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n708), .B1(new_n409), .B2(new_n413), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n413), .A2(new_n708), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n472), .B1(new_n818), .B2(new_n433), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n819), .B2(new_n777), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n710), .A2(new_n815), .A3(new_n777), .A4(new_n473), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT48), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n812), .B(new_n814), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n600), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n773), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n812), .A2(new_n814), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(KEYINPUT48), .A3(new_n821), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n829), .A3(new_n825), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n793), .B2(new_n794), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n754), .A2(KEYINPUT112), .A3(new_n760), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n792), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n796), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n804), .A2(new_n805), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n809), .A2(new_n833), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT118), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n690), .A2(new_n664), .A3(new_n713), .A4(new_n714), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n584), .B(new_n641), .C1(new_n362), .C2(new_n363), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n434), .A2(new_n845), .A3(new_n310), .A4(new_n637), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n631), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n717), .A2(new_n720), .A3(new_n724), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n649), .A2(new_n586), .ZN(new_n850));
  INV_X1    g664(.A(new_n640), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n631), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n658), .A2(new_n850), .A3(new_n713), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n643), .A2(new_n703), .A3(new_n665), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n526), .B1(new_n368), .B2(new_n366), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n580), .A2(new_n582), .A3(new_n824), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n568), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n568), .A3(KEYINPUT109), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n520), .A2(new_n682), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n580), .A2(new_n582), .A3(new_n860), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n699), .A2(new_n869), .A3(new_n632), .A4(new_n677), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n672), .A2(new_n675), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n849), .A2(new_n859), .A3(new_n866), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT53), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n875));
  OAI211_X1 g689(.A(new_n874), .B(KEYINPUT54), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n368), .A2(new_n366), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n567), .A3(new_n310), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n627), .A2(new_n631), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n677), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n871), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n699), .A3(new_n883), .A4(new_n869), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n864), .B2(new_n865), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n849), .A4(new_n859), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n809), .A2(new_n833), .A3(new_n891), .A4(new_n841), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n843), .A2(new_n876), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n813), .A2(new_n316), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n785), .A2(new_n566), .A3(new_n739), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n695), .B(KEYINPUT49), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n472), .A2(new_n584), .A3(new_n190), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n765), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(G75));
  NAND4_X1  g714(.A1(new_n877), .A2(new_n887), .A3(G902), .A4(new_n358), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n347), .A2(new_n352), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n350), .A2(new_n349), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n901), .B2(new_n902), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n316), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G51));
  XOR2_X1   g724(.A(new_n289), .B(KEYINPUT57), .Z(new_n911));
  AND3_X1   g725(.A1(new_n877), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT54), .B1(new_n877), .B2(new_n887), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n306), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n888), .A2(new_n308), .A3(new_n731), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n877), .A2(new_n887), .A3(G902), .A4(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n543), .A2(new_n560), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n919), .A2(KEYINPUT119), .A3(new_n920), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT119), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n909), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n595), .B(new_n927), .C1(new_n912), .C2(new_n913), .ZN(new_n928));
  INV_X1    g742(.A(new_n909), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n890), .B2(new_n876), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n595), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n877), .A2(new_n887), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n909), .B1(new_n936), .B2(new_n463), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n877), .A2(new_n887), .A3(new_n629), .A4(new_n935), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT61), .B1(new_n938), .B2(KEYINPUT120), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n937), .B(new_n938), .C1(KEYINPUT120), .C2(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  AOI21_X1  g757(.A(new_n316), .B1(new_n523), .B2(G224), .ZN(new_n944));
  INV_X1    g758(.A(new_n885), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n316), .ZN(new_n946));
  INV_X1    g760(.A(G898), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n903), .B1(new_n947), .B2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  MUX2_X1   g763(.A(new_n385), .B(new_n414), .S(KEYINPUT30), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n549), .A2(new_n553), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n717), .A2(new_n720), .A3(new_n724), .A4(new_n761), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n714), .B1(new_n743), .B2(new_n744), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n758), .A2(new_n578), .A3(new_n646), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT44), .B1(new_n746), .B2(new_n742), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n703), .A2(new_n643), .A3(new_n665), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n748), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n953), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n819), .A2(new_n736), .A3(new_n850), .ZN(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT127), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n959), .A2(new_n962), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n717), .A2(new_n720), .A3(new_n724), .A4(new_n761), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n964), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n316), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n968), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n952), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n952), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n434), .A2(new_n473), .A3(new_n714), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n867), .A2(KEYINPUT121), .A3(new_n600), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n310), .A3(new_n646), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT121), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n868), .B2(new_n824), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n979), .A2(KEYINPUT122), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n434), .A3(new_n473), .A4(new_n714), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n981), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n748), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n748), .A2(new_n985), .A3(new_n988), .A4(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n761), .ZN(new_n994));
  INV_X1    g808(.A(new_n660), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n960), .A3(KEYINPUT62), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n660), .B2(new_n958), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n993), .A2(new_n999), .A3(KEYINPUT124), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n978), .B1(new_n1004), .B2(new_n316), .ZN(new_n1005));
  OAI21_X1  g819(.A(G953), .B1(new_n280), .B2(new_n966), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n977), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1006), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n975), .B1(new_n974), .B2(new_n968), .ZN(new_n1009));
  AOI211_X1 g823(.A(KEYINPUT127), .B(new_n969), .C1(new_n973), .C2(new_n316), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n978), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1003), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT124), .B1(new_n993), .B2(new_n999), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n316), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n952), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1008), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1007), .A2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n945), .B2(new_n973), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n425), .A3(new_n430), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n431), .B1(new_n397), .B2(new_n398), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n874), .B(new_n1019), .C1(new_n873), .C2(new_n875), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1021), .B(new_n929), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1002), .A2(new_n885), .A3(new_n1003), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n430), .B1(new_n1025), .B2(new_n1019), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n1026), .B2(new_n391), .ZN(G57));
endmodule


