

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769;

  NAND2_X1 U372 ( .A1(n599), .A2(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U373 ( .A1(n711), .A2(n351), .ZN(n599) );
  AND2_X2 U374 ( .A1(n429), .A2(n427), .ZN(n426) );
  INV_X1 U375 ( .A(n625), .ZN(n680) );
  INV_X1 U376 ( .A(G953), .ZN(n760) );
  AND2_X1 U377 ( .A1(n635), .A2(n718), .ZN(n636) );
  AND2_X1 U378 ( .A1(n387), .A2(n386), .ZN(n349) );
  AND2_X2 U379 ( .A1(n664), .A2(n661), .ZN(n443) );
  NAND2_X2 U380 ( .A1(n587), .A2(n586), .ZN(n711) );
  XNOR2_X2 U381 ( .A(n584), .B(n583), .ZN(n587) );
  XNOR2_X2 U382 ( .A(n544), .B(n569), .ZN(n751) );
  XOR2_X2 U383 ( .A(G125), .B(G146), .Z(n519) );
  NOR2_X2 U384 ( .A1(n422), .A2(G953), .ZN(n421) );
  XNOR2_X2 U385 ( .A(n508), .B(n507), .ZN(n544) );
  XNOR2_X2 U386 ( .A(n554), .B(n505), .ZN(n508) );
  XNOR2_X2 U387 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n423) );
  XNOR2_X1 U388 ( .A(n590), .B(KEYINPUT32), .ZN(n351) );
  XNOR2_X1 U389 ( .A(n625), .B(n398), .ZN(n595) );
  INV_X1 U390 ( .A(KEYINPUT74), .ZN(n505) );
  INV_X1 U391 ( .A(G104), .ZN(n397) );
  AND2_X1 U392 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U393 ( .A1(n425), .A2(n466), .ZN(n424) );
  NAND2_X1 U394 ( .A1(n660), .A2(n358), .ZN(n664) );
  AND2_X1 U395 ( .A1(n390), .A2(n388), .ZN(n469) );
  XNOR2_X1 U396 ( .A(n591), .B(n402), .ZN(n418) );
  AND2_X1 U397 ( .A1(n389), .A2(n470), .ZN(n388) );
  NOR2_X2 U398 ( .A1(n589), .A2(n674), .ZN(n584) );
  BUF_X1 U399 ( .A(n575), .Z(n597) );
  NOR2_X1 U400 ( .A1(n640), .A2(n631), .ZN(n458) );
  AND2_X1 U401 ( .A1(n674), .A2(n477), .ZN(n596) );
  AND2_X1 U402 ( .A1(n613), .A2(n614), .ZN(n459) );
  NOR2_X1 U403 ( .A1(n549), .A2(n595), .ZN(n477) );
  AND2_X1 U404 ( .A1(n673), .A2(n612), .ZN(n613) );
  XNOR2_X1 U405 ( .A(n531), .B(n530), .ZN(n736) );
  XNOR2_X1 U406 ( .A(n465), .B(n464), .ZN(n745) );
  XNOR2_X1 U407 ( .A(n750), .B(n523), .ZN(n531) );
  XNOR2_X1 U408 ( .A(n357), .B(n478), .ZN(n539) );
  XNOR2_X1 U409 ( .A(n449), .B(G101), .ZN(n509) );
  XNOR2_X1 U410 ( .A(n397), .B(G110), .ZN(n510) );
  XOR2_X1 U411 ( .A(G119), .B(KEYINPUT3), .Z(n357) );
  INV_X1 U412 ( .A(G146), .ZN(n448) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n579) );
  XNOR2_X1 U414 ( .A(G107), .B(G122), .ZN(n481) );
  NOR2_X2 U415 ( .A1(n653), .A2(n764), .ZN(n657) );
  NAND2_X1 U416 ( .A1(n426), .A2(n424), .ZN(n431) );
  BUF_X1 U417 ( .A(n489), .Z(n350) );
  XNOR2_X1 U418 ( .A(n440), .B(n745), .ZN(n489) );
  XNOR2_X2 U419 ( .A(n614), .B(KEYINPUT1), .ZN(n674) );
  NOR2_X1 U420 ( .A1(n688), .A2(n671), .ZN(n476) );
  AND2_X1 U421 ( .A1(n416), .A2(n417), .ZN(n415) );
  XNOR2_X1 U422 ( .A(n351), .B(G119), .ZN(n765) );
  NOR2_X1 U423 ( .A1(n597), .A2(n537), .ZN(n538) );
  INV_X1 U424 ( .A(n669), .ZN(n352) );
  AND2_X1 U425 ( .A1(n598), .A2(n705), .ZN(n420) );
  NOR2_X2 U426 ( .A1(n489), .A2(n661), .ZN(n493) );
  NAND2_X2 U427 ( .A1(n643), .A2(n685), .ZN(n650) );
  XNOR2_X1 U428 ( .A(G469), .B(KEYINPUT75), .ZN(n513) );
  NOR2_X1 U429 ( .A1(n726), .A2(G902), .ZN(n514) );
  XNOR2_X1 U430 ( .A(n509), .B(n448), .ZN(n543) );
  NAND2_X1 U431 ( .A1(n690), .A2(n473), .ZN(n470) );
  NAND2_X1 U432 ( .A1(n471), .A2(n472), .ZN(n468) );
  NOR2_X1 U433 ( .A1(n707), .A2(KEYINPUT107), .ZN(n472) );
  INV_X1 U434 ( .A(G224), .ZN(n422) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n498) );
  INV_X1 U436 ( .A(KEYINPUT70), .ZN(n449) );
  XNOR2_X1 U437 ( .A(n622), .B(KEYINPUT38), .ZN(n686) );
  XNOR2_X1 U438 ( .A(n542), .B(n540), .ZN(n454) );
  XNOR2_X1 U439 ( .A(G113), .B(KEYINPUT76), .ZN(n478) );
  NAND2_X1 U440 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n751), .B(n436), .ZN(n726) );
  XNOR2_X1 U442 ( .A(n411), .B(n410), .ZN(n512) );
  XNOR2_X1 U443 ( .A(n511), .B(KEYINPUT97), .ZN(n410) );
  INV_X1 U444 ( .A(KEYINPUT89), .ZN(n444) );
  XNOR2_X1 U445 ( .A(n627), .B(n438), .ZN(n628) );
  XNOR2_X1 U446 ( .A(n439), .B(KEYINPUT113), .ZN(n438) );
  INV_X1 U447 ( .A(KEYINPUT121), .ZN(n435) );
  NAND2_X1 U448 ( .A1(n734), .A2(n395), .ZN(n394) );
  AND2_X1 U449 ( .A1(n662), .A2(G210), .ZN(n395) );
  AND2_X1 U450 ( .A1(n393), .A2(n407), .ZN(n392) );
  OR2_X1 U451 ( .A1(n662), .A2(G210), .ZN(n393) );
  INV_X1 U452 ( .A(KEYINPUT66), .ZN(n402) );
  NOR2_X1 U453 ( .A1(n768), .A2(n767), .ZN(n401) );
  XNOR2_X1 U454 ( .A(G122), .B(G113), .ZN(n562) );
  XOR2_X1 U455 ( .A(G143), .B(KEYINPUT12), .Z(n563) );
  XNOR2_X1 U456 ( .A(G131), .B(G140), .ZN(n569) );
  XNOR2_X1 U457 ( .A(n543), .B(n510), .ZN(n411) );
  XNOR2_X1 U458 ( .A(G902), .B(KEYINPUT15), .ZN(n515) );
  XNOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT94), .ZN(n437) );
  NOR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n490) );
  INV_X1 U461 ( .A(KEYINPUT28), .ZN(n439) );
  XNOR2_X1 U462 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n501) );
  INV_X1 U463 ( .A(KEYINPUT6), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n604), .B(KEYINPUT45), .ZN(n475) );
  XNOR2_X1 U465 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n524) );
  XNOR2_X1 U466 ( .A(G110), .B(G128), .ZN(n521) );
  XOR2_X1 U467 ( .A(G137), .B(G140), .Z(n522) );
  INV_X1 U468 ( .A(G134), .ZN(n503) );
  XNOR2_X1 U469 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n552) );
  XOR2_X1 U470 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n527) );
  INV_X1 U471 ( .A(n686), .ZN(n631) );
  INV_X1 U472 ( .A(n641), .ZN(n446) );
  INV_X1 U473 ( .A(KEYINPUT109), .ZN(n583) );
  XNOR2_X1 U474 ( .A(n574), .B(n433), .ZN(n576) );
  XNOR2_X1 U475 ( .A(n573), .B(G475), .ZN(n433) );
  XNOR2_X1 U476 ( .A(n455), .B(n453), .ZN(n545) );
  XNOR2_X1 U477 ( .A(n454), .B(n541), .ZN(n453) );
  XNOR2_X1 U478 ( .A(n543), .B(n456), .ZN(n455) );
  XNOR2_X1 U479 ( .A(n482), .B(n479), .ZN(n464) );
  NAND2_X1 U480 ( .A1(n381), .A2(n367), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n734), .A2(n382), .ZN(n381) );
  OR2_X1 U482 ( .A1(n729), .A2(G475), .ZN(n380) );
  INV_X1 U483 ( .A(n376), .ZN(n375) );
  NAND2_X1 U484 ( .A1(n379), .A2(n406), .ZN(n373) );
  AND2_X1 U485 ( .A1(n376), .A2(n730), .ZN(n370) );
  NOR2_X1 U486 ( .A1(n428), .A2(G953), .ZN(n427) );
  NOR2_X1 U487 ( .A1(n353), .A2(KEYINPUT119), .ZN(n428) );
  NAND2_X2 U488 ( .A1(n349), .A2(n383), .ZN(n721) );
  NOR2_X1 U489 ( .A1(n669), .A2(n364), .ZN(n384) );
  NOR2_X1 U490 ( .A1(n633), .A2(n432), .ZN(n716) );
  XNOR2_X1 U491 ( .A(n731), .B(n434), .ZN(n733) );
  XNOR2_X1 U492 ( .A(n732), .B(n435), .ZN(n434) );
  AND2_X1 U493 ( .A1(n403), .A2(n407), .ZN(G54) );
  XNOR2_X1 U494 ( .A(n405), .B(n404), .ZN(n403) );
  XNOR2_X1 U495 ( .A(n726), .B(n368), .ZN(n404) );
  NOR2_X1 U496 ( .A1(n396), .A2(n391), .ZN(n663) );
  NOR2_X1 U497 ( .A1(n734), .A2(n662), .ZN(n396) );
  NOR2_X1 U498 ( .A1(n703), .A2(n362), .ZN(n353) );
  AND2_X1 U499 ( .A1(n474), .A2(KEYINPUT107), .ZN(n354) );
  AND2_X1 U500 ( .A1(n674), .A2(n361), .ZN(n355) );
  XOR2_X1 U501 ( .A(n492), .B(n491), .Z(n356) );
  NOR2_X1 U502 ( .A1(n659), .A2(n658), .ZN(n358) );
  XOR2_X1 U503 ( .A(n506), .B(n437), .Z(n359) );
  INV_X1 U504 ( .A(n690), .ZN(n474) );
  NOR2_X1 U505 ( .A1(n669), .A2(n668), .ZN(n360) );
  AND2_X1 U506 ( .A1(n670), .A2(n595), .ZN(n361) );
  AND2_X1 U507 ( .A1(n683), .A2(n694), .ZN(n362) );
  AND2_X1 U508 ( .A1(n353), .A2(KEYINPUT119), .ZN(n363) );
  INV_X1 U509 ( .A(KEYINPUT107), .ZN(n473) );
  XOR2_X1 U510 ( .A(n551), .B(KEYINPUT31), .Z(n364) );
  XOR2_X1 U511 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n365) );
  XOR2_X1 U512 ( .A(n704), .B(KEYINPUT62), .Z(n366) );
  AND2_X1 U513 ( .A1(n380), .A2(n407), .ZN(n367) );
  INV_X1 U514 ( .A(KEYINPUT92), .ZN(n447) );
  NOR2_X1 U515 ( .A1(G952), .A2(n760), .ZN(n738) );
  INV_X1 U516 ( .A(n738), .ZN(n407) );
  XNOR2_X1 U517 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n368) );
  INV_X1 U518 ( .A(n730), .ZN(n406) );
  INV_X1 U519 ( .A(KEYINPUT119), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n418), .A2(n447), .ZN(n413) );
  NAND2_X1 U521 ( .A1(n372), .A2(n369), .ZN(G60) );
  NAND2_X1 U522 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U523 ( .A(n379), .ZN(n371) );
  NAND2_X1 U524 ( .A1(n375), .A2(n406), .ZN(n374) );
  INV_X1 U525 ( .A(n729), .ZN(n377) );
  INV_X1 U526 ( .A(n734), .ZN(n378) );
  AND2_X1 U527 ( .A1(n729), .A2(G475), .ZN(n382) );
  NAND2_X1 U528 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U529 ( .A(n550), .ZN(n385) );
  NAND2_X1 U530 ( .A1(n669), .A2(n364), .ZN(n386) );
  NAND2_X1 U531 ( .A1(n550), .A2(n364), .ZN(n387) );
  NAND2_X1 U532 ( .A1(n721), .A2(n354), .ZN(n389) );
  NAND2_X1 U533 ( .A1(n707), .A2(n354), .ZN(n390) );
  XNOR2_X2 U534 ( .A(n548), .B(KEYINPUT101), .ZN(n707) );
  NAND2_X1 U535 ( .A1(n394), .A2(n392), .ZN(n391) );
  AND2_X4 U536 ( .A1(n445), .A2(n443), .ZN(n734) );
  NAND2_X1 U537 ( .A1(n414), .A2(n413), .ZN(n412) );
  XNOR2_X1 U538 ( .A(n510), .B(KEYINPUT16), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n408), .B(KEYINPUT35), .ZN(n601) );
  NOR2_X1 U540 ( .A1(n704), .A2(G902), .ZN(n546) );
  XNOR2_X1 U541 ( .A(n399), .B(n365), .ZN(n409) );
  NOR2_X1 U542 ( .A1(n667), .A2(n597), .ZN(n399) );
  NOR2_X1 U543 ( .A1(n666), .A2(n633), .ZN(n634) );
  XNOR2_X1 U544 ( .A(n632), .B(KEYINPUT41), .ZN(n666) );
  XNOR2_X1 U545 ( .A(n400), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n423), .B(n421), .ZN(n400) );
  XNOR2_X1 U547 ( .A(n401), .B(KEYINPUT46), .ZN(n646) );
  XNOR2_X1 U548 ( .A(n480), .B(n539), .ZN(n465) );
  XNOR2_X1 U549 ( .A(n431), .B(n430), .ZN(G75) );
  NAND2_X1 U550 ( .A1(n734), .A2(G469), .ZN(n405) );
  NAND2_X1 U551 ( .A1(n409), .A2(n446), .ZN(n408) );
  NAND2_X1 U552 ( .A1(n415), .A2(n412), .ZN(n442) );
  INV_X1 U553 ( .A(n419), .ZN(n414) );
  NAND2_X1 U554 ( .A1(n418), .A2(n447), .ZN(n416) );
  NAND2_X1 U555 ( .A1(n419), .A2(n447), .ZN(n417) );
  NAND2_X1 U556 ( .A1(n582), .A2(n420), .ZN(n419) );
  INV_X1 U557 ( .A(n467), .ZN(n425) );
  NAND2_X1 U558 ( .A1(n467), .A2(n363), .ZN(n429) );
  INV_X1 U559 ( .A(KEYINPUT53), .ZN(n430) );
  XNOR2_X1 U560 ( .A(n450), .B(KEYINPUT48), .ZN(n653) );
  INV_X1 U561 ( .A(n539), .ZN(n456) );
  NOR2_X1 U562 ( .A1(n723), .A2(n452), .ZN(n451) );
  XNOR2_X1 U563 ( .A(n512), .B(G107), .ZN(n436) );
  XNOR2_X2 U564 ( .A(n654), .B(KEYINPUT90), .ZN(n753) );
  BUF_X1 U565 ( .A(n629), .Z(n432) );
  XNOR2_X1 U566 ( .A(n486), .B(n359), .ZN(n440) );
  NAND2_X1 U567 ( .A1(n646), .A2(n451), .ZN(n450) );
  NAND2_X1 U568 ( .A1(n645), .A2(n647), .ZN(n452) );
  NOR2_X1 U569 ( .A1(n739), .A2(n753), .ZN(n655) );
  XNOR2_X2 U570 ( .A(n441), .B(n475), .ZN(n739) );
  NOR2_X2 U571 ( .A1(n629), .A2(n500), .ZN(n502) );
  NAND2_X1 U572 ( .A1(n442), .A2(n603), .ZN(n441) );
  XNOR2_X1 U573 ( .A(n445), .B(n444), .ZN(n665) );
  OR2_X2 U574 ( .A1(n655), .A2(KEYINPUT2), .ZN(n445) );
  INV_X1 U575 ( .A(n674), .ZN(n669) );
  XNOR2_X2 U576 ( .A(n514), .B(n513), .ZN(n614) );
  XNOR2_X1 U577 ( .A(n458), .B(n457), .ZN(n635) );
  INV_X1 U578 ( .A(KEYINPUT39), .ZN(n457) );
  NAND2_X1 U579 ( .A1(n460), .A2(n459), .ZN(n640) );
  XNOR2_X1 U580 ( .A(n605), .B(n606), .ZN(n460) );
  XNOR2_X1 U581 ( .A(n461), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U582 ( .A1(n462), .A2(n407), .ZN(n461) );
  XNOR2_X1 U583 ( .A(n463), .B(n366), .ZN(n462) );
  NAND2_X1 U584 ( .A1(n734), .A2(G472), .ZN(n463) );
  XNOR2_X2 U585 ( .A(n520), .B(KEYINPUT10), .ZN(n750) );
  INV_X1 U586 ( .A(n643), .ZN(n622) );
  XNOR2_X2 U587 ( .A(n650), .B(n495), .ZN(n629) );
  XNOR2_X2 U588 ( .A(n493), .B(n356), .ZN(n643) );
  NAND2_X1 U589 ( .A1(n665), .A2(n664), .ZN(n467) );
  NAND2_X1 U590 ( .A1(n469), .A2(n468), .ZN(n582) );
  INV_X1 U591 ( .A(n721), .ZN(n471) );
  INV_X1 U592 ( .A(n504), .ZN(n483) );
  XNOR2_X1 U593 ( .A(n545), .B(n544), .ZN(n704) );
  INV_X1 U594 ( .A(KEYINPUT102), .ZN(n551) );
  XNOR2_X1 U595 ( .A(n728), .B(n727), .ZN(n729) );
  INV_X1 U596 ( .A(n670), .ZN(n585) );
  NOR2_X1 U597 ( .A1(n680), .A2(n585), .ZN(n586) );
  XOR2_X1 U598 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n488) );
  XOR2_X1 U599 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n479) );
  XNOR2_X1 U600 ( .A(n481), .B(G116), .ZN(n559) );
  INV_X1 U601 ( .A(n559), .ZN(n482) );
  XOR2_X1 U602 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n506) );
  XOR2_X2 U603 ( .A(G143), .B(G128), .Z(n504) );
  XNOR2_X1 U604 ( .A(n519), .B(n509), .ZN(n484) );
  XNOR2_X1 U605 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U606 ( .A(n350), .B(KEYINPUT93), .ZN(n487) );
  XNOR2_X1 U607 ( .A(n488), .B(n487), .ZN(n662) );
  XNOR2_X1 U608 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n495) );
  INV_X1 U609 ( .A(n515), .ZN(n661) );
  XOR2_X1 U610 ( .A(KEYINPUT87), .B(KEYINPUT95), .Z(n492) );
  XNOR2_X1 U611 ( .A(n490), .B(KEYINPUT81), .ZN(n494) );
  NAND2_X1 U612 ( .A1(G210), .A2(n494), .ZN(n491) );
  NAND2_X1 U613 ( .A1(G214), .A2(n494), .ZN(n685) );
  NOR2_X1 U614 ( .A1(G898), .A2(n760), .ZN(n496) );
  XNOR2_X1 U615 ( .A(KEYINPUT96), .B(n496), .ZN(n746) );
  NAND2_X1 U616 ( .A1(n746), .A2(G902), .ZN(n497) );
  NAND2_X1 U617 ( .A1(G952), .A2(n760), .ZN(n608) );
  AND2_X1 U618 ( .A1(n497), .A2(n608), .ZN(n499) );
  XNOR2_X1 U619 ( .A(n498), .B(KEYINPUT14), .ZN(n610) );
  INV_X1 U620 ( .A(n610), .ZN(n702) );
  OR2_X1 U621 ( .A1(n499), .A2(n702), .ZN(n500) );
  XNOR2_X1 U622 ( .A(n502), .B(n501), .ZN(n575) );
  XNOR2_X2 U623 ( .A(n504), .B(n503), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n506), .B(G137), .ZN(n507) );
  NAND2_X1 U625 ( .A1(G227), .A2(n760), .ZN(n511) );
  XOR2_X1 U626 ( .A(KEYINPUT21), .B(KEYINPUT99), .Z(n518) );
  NAND2_X1 U627 ( .A1(G234), .A2(n515), .ZN(n516) );
  XNOR2_X1 U628 ( .A(KEYINPUT20), .B(n516), .ZN(n532) );
  NAND2_X1 U629 ( .A1(n532), .A2(G221), .ZN(n517) );
  XNOR2_X1 U630 ( .A(n518), .B(n517), .ZN(n671) );
  XNOR2_X1 U631 ( .A(n519), .B(KEYINPUT73), .ZN(n520) );
  XNOR2_X1 U632 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U633 ( .A(n524), .B(KEYINPUT98), .ZN(n525) );
  XOR2_X1 U634 ( .A(G119), .B(n525), .Z(n529) );
  NAND2_X1 U635 ( .A1(G234), .A2(n760), .ZN(n526) );
  XNOR2_X1 U636 ( .A(n527), .B(n526), .ZN(n555) );
  NAND2_X1 U637 ( .A1(G221), .A2(n555), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U639 ( .A1(n736), .A2(G902), .ZN(n536) );
  XOR2_X1 U640 ( .A(KEYINPUT25), .B(KEYINPUT84), .Z(n534) );
  NAND2_X1 U641 ( .A1(n532), .A2(G217), .ZN(n533) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X2 U643 ( .A(n536), .B(n535), .ZN(n670) );
  NOR2_X2 U644 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U645 ( .A1(n614), .A2(n673), .ZN(n537) );
  XNOR2_X1 U646 ( .A(n538), .B(KEYINPUT100), .ZN(n547) );
  XOR2_X1 U647 ( .A(KEYINPUT82), .B(KEYINPUT5), .Z(n541) );
  XNOR2_X1 U648 ( .A(G116), .B(G131), .ZN(n540) );
  NOR2_X1 U649 ( .A1(G953), .A2(G237), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n565), .A2(G210), .ZN(n542) );
  XNOR2_X2 U651 ( .A(n546), .B(G472), .ZN(n625) );
  NAND2_X1 U652 ( .A1(n547), .A2(n625), .ZN(n548) );
  INV_X1 U653 ( .A(n673), .ZN(n549) );
  OR2_X1 U654 ( .A1(n625), .A2(n549), .ZN(n668) );
  OR2_X1 U655 ( .A1(n597), .A2(n668), .ZN(n550) );
  XNOR2_X1 U656 ( .A(n552), .B(KEYINPUT105), .ZN(n553) );
  XOR2_X1 U657 ( .A(n554), .B(n553), .Z(n557) );
  NAND2_X1 U658 ( .A1(G217), .A2(n555), .ZN(n556) );
  XNOR2_X1 U659 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U660 ( .A(n559), .B(n558), .ZN(n732) );
  NOR2_X1 U661 ( .A1(G902), .A2(n732), .ZN(n561) );
  XNOR2_X1 U662 ( .A(KEYINPUT106), .B(G478), .ZN(n560) );
  XNOR2_X1 U663 ( .A(n561), .B(n560), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U665 ( .A(n750), .B(n564), .ZN(n572) );
  XOR2_X1 U666 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n567) );
  NAND2_X1 U667 ( .A1(n565), .A2(G214), .ZN(n566) );
  XNOR2_X1 U668 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U669 ( .A(G104), .B(n568), .ZN(n570) );
  XNOR2_X1 U670 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n572), .B(n571), .ZN(n728) );
  NOR2_X1 U672 ( .A1(G902), .A2(n728), .ZN(n574) );
  XNOR2_X1 U673 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n573) );
  NAND2_X1 U674 ( .A1(n593), .A2(n576), .ZN(n617) );
  INV_X1 U675 ( .A(n617), .ZN(n718) );
  NOR2_X1 U676 ( .A1(n593), .A2(n576), .ZN(n720) );
  NOR2_X1 U677 ( .A1(n718), .A2(n720), .ZN(n690) );
  INV_X1 U678 ( .A(n575), .ZN(n578) );
  INV_X1 U679 ( .A(n576), .ZN(n592) );
  NAND2_X1 U680 ( .A1(n592), .A2(n593), .ZN(n577) );
  XNOR2_X1 U681 ( .A(n577), .B(KEYINPUT108), .ZN(n688) );
  NAND2_X1 U682 ( .A1(n578), .A2(n476), .ZN(n580) );
  XNOR2_X1 U683 ( .A(n580), .B(n579), .ZN(n589) );
  INV_X1 U684 ( .A(n595), .ZN(n619) );
  NOR2_X1 U685 ( .A1(n619), .A2(n670), .ZN(n581) );
  NAND2_X1 U686 ( .A1(n584), .A2(n581), .ZN(n705) );
  XOR2_X1 U687 ( .A(KEYINPUT86), .B(n355), .Z(n588) );
  OR2_X1 U688 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U689 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U690 ( .A(KEYINPUT110), .B(n594), .Z(n641) );
  XNOR2_X1 U691 ( .A(n596), .B(KEYINPUT33), .ZN(n667) );
  NAND2_X1 U692 ( .A1(n601), .A2(KEYINPUT44), .ZN(n598) );
  BUF_X1 U693 ( .A(n599), .Z(n600) );
  NOR2_X1 U694 ( .A1(KEYINPUT44), .A2(n600), .ZN(n602) );
  INV_X1 U695 ( .A(n601), .ZN(n766) );
  NAND2_X1 U696 ( .A1(n602), .A2(n766), .ZN(n603) );
  XNOR2_X1 U697 ( .A(KEYINPUT91), .B(KEYINPUT64), .ZN(n604) );
  XOR2_X1 U698 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n606) );
  NAND2_X1 U699 ( .A1(n680), .A2(n685), .ZN(n605) );
  NOR2_X1 U700 ( .A1(G900), .A2(n760), .ZN(n607) );
  NAND2_X1 U701 ( .A1(n607), .A2(G902), .ZN(n609) );
  NAND2_X1 U702 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U703 ( .A1(n611), .A2(n610), .ZN(n615) );
  INV_X1 U704 ( .A(n615), .ZN(n612) );
  NAND2_X1 U705 ( .A1(n635), .A2(n720), .ZN(n725) );
  NOR2_X1 U706 ( .A1(n671), .A2(n615), .ZN(n616) );
  NAND2_X1 U707 ( .A1(n616), .A2(n670), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n626), .A2(n617), .ZN(n618) );
  NAND2_X1 U709 ( .A1(n619), .A2(n618), .ZN(n648) );
  NOR2_X1 U710 ( .A1(n352), .A2(n648), .ZN(n620) );
  NAND2_X1 U711 ( .A1(n620), .A2(n685), .ZN(n621) );
  XNOR2_X1 U712 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U714 ( .A(KEYINPUT111), .B(n624), .ZN(n764) );
  NOR2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U716 ( .A1(n628), .A2(n614), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n474), .A2(n716), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n630), .A2(KEYINPUT47), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n686), .A2(n685), .ZN(n689) );
  NOR2_X1 U720 ( .A1(n689), .A2(n688), .ZN(n632) );
  XNOR2_X1 U721 ( .A(n634), .B(KEYINPUT42), .ZN(n768) );
  XNOR2_X1 U722 ( .A(n636), .B(KEYINPUT40), .ZN(n767) );
  XOR2_X1 U723 ( .A(KEYINPUT47), .B(KEYINPUT71), .Z(n637) );
  NOR2_X1 U724 ( .A1(n690), .A2(n637), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT80), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n639), .A2(n716), .ZN(n644) );
  NOR2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n715) );
  AND2_X1 U729 ( .A1(n644), .A2(n715), .ZN(n645) );
  XNOR2_X1 U730 ( .A(KEYINPUT114), .B(n648), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT36), .B(n651), .Z(n652) );
  NOR2_X1 U733 ( .A1(n669), .A2(n652), .ZN(n723) );
  NAND2_X1 U734 ( .A1(n725), .A2(n657), .ZN(n654) );
  INV_X1 U735 ( .A(n739), .ZN(n660) );
  NAND2_X1 U736 ( .A1(KEYINPUT2), .A2(n725), .ZN(n656) );
  XNOR2_X1 U737 ( .A(KEYINPUT88), .B(n656), .ZN(n659) );
  INV_X1 U738 ( .A(n657), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U740 ( .A(n666), .ZN(n683) );
  INV_X1 U741 ( .A(n667), .ZN(n694) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(n672), .Z(n678) );
  XNOR2_X1 U744 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n352), .A2(n673), .ZN(n675) );
  XOR2_X1 U746 ( .A(n676), .B(n675), .Z(n677) );
  NAND2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n360), .A2(n681), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT51), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n697) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(KEYINPUT117), .B(n693), .ZN(n695) );
  NAND2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n699), .B(KEYINPUT118), .ZN(n700) );
  NAND2_X1 U761 ( .A1(n700), .A2(G952), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U763 ( .A(G101), .B(n705), .ZN(G3) );
  NAND2_X1 U764 ( .A1(n707), .A2(n718), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n706), .B(G104), .ZN(G6) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U767 ( .A1(n707), .A2(n720), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U769 ( .A(G107), .B(n710), .ZN(G9) );
  XNOR2_X1 U770 ( .A(n711), .B(G110), .ZN(G12) );
  XOR2_X1 U771 ( .A(G128), .B(KEYINPUT29), .Z(n713) );
  NAND2_X1 U772 ( .A1(n716), .A2(n720), .ZN(n712) );
  XNOR2_X1 U773 ( .A(n713), .B(n712), .ZN(G30) );
  XOR2_X1 U774 ( .A(G143), .B(KEYINPUT115), .Z(n714) );
  XNOR2_X1 U775 ( .A(n715), .B(n714), .ZN(G45) );
  NAND2_X1 U776 ( .A1(n716), .A2(n718), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n717), .B(G146), .ZN(G48) );
  NAND2_X1 U778 ( .A1(n721), .A2(n718), .ZN(n719) );
  XNOR2_X1 U779 ( .A(n719), .B(G113), .ZN(G15) );
  NAND2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n722), .B(G116), .ZN(G18) );
  XNOR2_X1 U782 ( .A(G125), .B(n723), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U784 ( .A(G134), .B(n725), .ZN(G36) );
  XNOR2_X1 U785 ( .A(KEYINPUT59), .B(KEYINPUT120), .ZN(n727) );
  XNOR2_X1 U786 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n730) );
  NAND2_X1 U787 ( .A1(n734), .A2(G478), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n738), .A2(n733), .ZN(G63) );
  NAND2_X1 U789 ( .A1(G217), .A2(n734), .ZN(n735) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n738), .A2(n737), .ZN(G66) );
  OR2_X1 U792 ( .A1(G953), .A2(n739), .ZN(n743) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n740) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n740), .ZN(n741) );
  NAND2_X1 U795 ( .A1(n741), .A2(G898), .ZN(n742) );
  NAND2_X1 U796 ( .A1(n743), .A2(n742), .ZN(n749) );
  XOR2_X1 U797 ( .A(G101), .B(KEYINPUT122), .Z(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(G69) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(n756) );
  INV_X1 U802 ( .A(n756), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U804 ( .A1(G953), .A2(n754), .ZN(n755) );
  XNOR2_X1 U805 ( .A(KEYINPUT123), .B(n755), .ZN(n763) );
  XNOR2_X1 U806 ( .A(G227), .B(n756), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n757), .A2(G900), .ZN(n758) );
  XOR2_X1 U808 ( .A(KEYINPUT124), .B(n758), .Z(n759) );
  NOR2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U810 ( .A(KEYINPUT125), .B(n761), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U812 ( .A(G140), .B(n764), .Z(G42) );
  XNOR2_X1 U813 ( .A(n765), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U814 ( .A(G122), .B(n766), .ZN(G24) );
  XOR2_X1 U815 ( .A(G131), .B(n767), .Z(G33) );
  XNOR2_X1 U816 ( .A(G137), .B(KEYINPUT127), .ZN(n769) );
  XNOR2_X1 U817 ( .A(n769), .B(n768), .ZN(G39) );
endmodule

