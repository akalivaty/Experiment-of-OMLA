//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR4_X1   g017(.A1(KEYINPUT90), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(new_n213), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n215), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT91), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(new_n215), .C1(new_n219), .C2(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n210), .ZN(new_n227));
  INV_X1    g026(.A(new_n209), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n218), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(KEYINPUT93), .C1(G1gat), .C2(new_n230), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT92), .B1(new_n229), .B2(KEYINPUT17), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n223), .A2(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n209), .B1(new_n240), .B2(new_n226), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n218), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n233), .B(G8gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(KEYINPUT17), .B2(new_n229), .ZN(new_n245));
  AOI211_X1 g044(.A(new_n204), .B(new_n236), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n202), .B1(new_n246), .B2(KEYINPUT18), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT11), .B(G169gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n215), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n214), .A2(KEYINPUT90), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n220), .A3(new_n213), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n210), .B1(new_n257), .B2(new_n225), .ZN(new_n258));
  INV_X1    g057(.A(new_n226), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n228), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n217), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n229), .A2(new_n235), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n203), .B(KEYINPUT13), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n246), .B2(KEYINPUT18), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n243), .A2(new_n245), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n247), .B(new_n253), .C1(new_n267), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n203), .A3(new_n262), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT18), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n272), .A2(new_n273), .B1(new_n264), .B2(new_n265), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT94), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n274), .B(new_n269), .C1(new_n275), .C2(new_n252), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT73), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(KEYINPUT26), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(KEYINPUT28), .A3(new_n290), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n290), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n287), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT23), .B1(new_n282), .B2(KEYINPUT65), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n296), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(new_n301), .B2(new_n297), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n295), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n281), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n314), .B2(new_n279), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT72), .B(G218gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT22), .B1(new_n317), .B2(G211gat), .ZN(new_n318));
  XOR2_X1   g117(.A(G197gat), .B(G204gat), .Z(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n318), .B2(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n314), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n280), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n279), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT74), .ZN(new_n332));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT30), .ZN(new_n336));
  OR3_X1    g135(.A1(new_n335), .A2(KEYINPUT76), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n334), .B(KEYINPUT75), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n326), .B2(new_n330), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n335), .B1(new_n339), .B2(new_n336), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n335), .B2(new_n336), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  INV_X1    g150(.A(G127gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT67), .B(G113gat), .Z(new_n355));
  OAI211_X1 g154(.A(new_n350), .B(new_n345), .C1(new_n355), .C2(new_n349), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n311), .A2(new_n303), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n358), .A2(new_n296), .B1(new_n311), .B2(new_n312), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n359), .B2(new_n295), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n356), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n314), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n344), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT68), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n369), .B1(new_n375), .B2(KEYINPUT69), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(KEYINPUT69), .B2(new_n375), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT32), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n365), .B2(new_n367), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n364), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT71), .B1(new_n382), .B2(KEYINPUT34), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n366), .B1(new_n360), .B2(new_n362), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT34), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n384), .B2(new_n386), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n381), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n392), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n374), .B1(new_n368), .B2(new_n370), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  INV_X1    g198(.A(G155gat), .ZN(new_n400));
  INV_X1    g199(.A(G162gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G141gat), .B(G148gat), .ZN(new_n406));
  OAI221_X1 g205(.A(new_n405), .B1(new_n403), .B2(new_n404), .C1(KEYINPUT2), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G148gat), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT78), .B1(new_n408), .B2(G141gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  INV_X1    g209(.A(G141gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(G148gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(G141gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT79), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT80), .B(G155gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT2), .B1(new_n416), .B2(new_n401), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n409), .A2(new_n412), .A3(new_n418), .A4(new_n413), .ZN(new_n419));
  XNOR2_X1  g218(.A(G155gat), .B(G162gat), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(new_n417), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n407), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n324), .A2(new_n399), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n421), .A3(new_n424), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n324), .B1(new_n428), .B2(new_n399), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n398), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(KEYINPUT3), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n423), .A2(G228gat), .A3(new_n432), .A4(G233gat), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT86), .B1(new_n428), .B2(new_n399), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n324), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(KEYINPUT86), .A3(new_n399), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(G22gat), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n435), .A2(new_n436), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n439), .B(new_n430), .C1(new_n440), .C2(new_n433), .ZN(new_n441));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT31), .B(G50gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND4_X1  g243(.A1(new_n438), .A2(new_n441), .A3(KEYINPUT87), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n441), .A3(KEYINPUT87), .ZN(new_n446));
  INV_X1    g245(.A(new_n444), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT87), .B1(new_n438), .B2(new_n441), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n397), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT0), .ZN(new_n453));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n357), .A2(new_n421), .A3(new_n407), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n407), .A2(new_n421), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n357), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n432), .A2(new_n428), .A3(new_n361), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n465), .A2(new_n464), .A3(new_n460), .A4(new_n462), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n422), .A2(new_n361), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  INV_X1    g269(.A(new_n464), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n457), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT83), .B1(new_n468), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n456), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT84), .B(new_n456), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(new_n482), .B2(new_n455), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT6), .B(new_n456), .C1(new_n474), .C2(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n343), .B(new_n451), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  NOR4_X1   g288(.A1(new_n397), .A2(new_n450), .A3(KEYINPUT35), .A4(new_n342), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(KEYINPUT88), .B(new_n456), .C1(new_n474), .C2(new_n475), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n483), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n393), .B2(new_n396), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n393), .A2(new_n396), .A3(new_n498), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n455), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT39), .B1(new_n470), .B2(new_n471), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT40), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n456), .B1(new_n503), .B2(new_n504), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(new_n511), .C1(new_n503), .C2(new_n507), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n342), .A2(new_n513), .A3(new_n492), .A4(new_n493), .ZN(new_n514));
  INV_X1    g313(.A(new_n450), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n326), .A2(new_n518), .A3(new_n330), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n316), .A2(new_n324), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n328), .A2(new_n325), .A3(new_n329), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT37), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n338), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n335), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n326), .A2(new_n330), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT37), .ZN(new_n528));
  INV_X1    g327(.A(new_n334), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n519), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n494), .A3(new_n485), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n502), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n343), .B1(new_n486), .B2(new_n487), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n450), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n278), .B1(new_n497), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G134gat), .B(G162gat), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(KEYINPUT41), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g343(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(G85gat), .A3(G92gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(new_n547), .A3(new_n551), .A4(new_n554), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n261), .B2(new_n239), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n237), .B2(new_n242), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n540), .A2(KEYINPUT41), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n229), .B2(new_n561), .ZN(new_n565));
  OAI21_X1  g364(.A(G190gat), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n229), .B2(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n243), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n565), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n290), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G218gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT99), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n570), .A3(G218gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n542), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n290), .B1(new_n568), .B2(new_n569), .ZN(new_n576));
  AOI211_X1 g375(.A(G190gat), .B(new_n565), .C1(new_n243), .C2(new_n567), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n574), .A3(new_n579), .A4(new_n542), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n539), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT96), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT97), .ZN(new_n592));
  NAND2_X1  g391(.A1(G57gat), .A2(G64gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT95), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(G57gat), .A2(G64gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n593), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n590), .A2(new_n592), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(KEYINPUT9), .A3(new_n593), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n585), .A3(new_n583), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT21), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n352), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n596), .A2(new_n599), .A3(new_n586), .A4(new_n589), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n591), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n602), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(KEYINPUT98), .B(new_n602), .C1(new_n607), .C2(new_n609), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT21), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n235), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n606), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G155gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n578), .A2(new_n579), .A3(new_n574), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n541), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n538), .A3(new_n580), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  INV_X1    g426(.A(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n600), .A2(new_n602), .A3(new_n557), .A4(new_n559), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n560), .A2(new_n610), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT10), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n557), .B2(new_n559), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n612), .A2(new_n613), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n630), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n631), .A2(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n629), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n639), .A3(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n582), .A2(new_n623), .A3(new_n626), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n537), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n486), .A2(new_n487), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(G1gat), .Z(G1324gat));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND4_X1  g455(.A1(new_n537), .A2(new_n342), .A3(new_n650), .A4(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G8gat), .B1(new_n651), .B2(new_n343), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n657), .ZN(new_n659));
  MUX2_X1   g458(.A(new_n657), .B(new_n659), .S(KEYINPUT42), .Z(G1325gat));
  AND3_X1   g459(.A1(new_n393), .A2(new_n396), .A3(new_n498), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n499), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n651), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n397), .A2(G15gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n651), .B2(new_n664), .ZN(G1326gat));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n651), .B2(new_n515), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n537), .A2(KEYINPUT102), .A3(new_n450), .A4(new_n650), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n582), .A2(new_n626), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n531), .A2(new_n494), .A3(new_n485), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n662), .B1(new_n673), .B2(new_n516), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n534), .B2(new_n450), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n488), .A2(KEYINPUT35), .B1(new_n495), .B2(new_n490), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(KEYINPUT44), .B(new_n672), .C1(new_n675), .C2(new_n676), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n623), .A2(new_n647), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n277), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n271), .A2(new_n276), .A3(KEYINPUT103), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n679), .A2(new_n652), .A3(new_n680), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G29gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n497), .A2(new_n536), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n681), .A2(new_n672), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n277), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n653), .A2(G29gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT45), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n537), .A2(new_n695), .A3(new_n690), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n688), .A2(new_n697), .A3(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n691), .A2(G36gat), .A3(new_n343), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n679), .A2(new_n680), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n705), .A2(new_n342), .A3(new_n686), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n213), .B2(new_n706), .ZN(G1329gat));
  OR3_X1    g506(.A1(new_n691), .A2(G43gat), .A3(new_n397), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT47), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n679), .A2(new_n502), .A3(new_n680), .A4(new_n686), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n708), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n712), .B(new_n708), .C1(new_n709), .C2(KEYINPUT47), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  OR3_X1    g515(.A1(new_n691), .A2(G50gat), .A3(new_n515), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n717), .A2(KEYINPUT48), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n679), .A2(new_n450), .A3(new_n680), .A4(new_n686), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G50gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1331gat));
  INV_X1    g528(.A(new_n623), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n672), .A2(new_n685), .A3(new_n730), .A4(new_n648), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n689), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n652), .A2(KEYINPUT107), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n652), .A2(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n738));
  INV_X1    g537(.A(G64gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n732), .B(new_n342), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1333gat));
  XOR2_X1   g541(.A(new_n397), .B(KEYINPUT109), .Z(new_n743));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(G71gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n689), .A2(G71gat), .A3(new_n502), .A4(new_n731), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT50), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n746), .B(new_n752), .C1(new_n748), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n732), .A2(new_n450), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n685), .A2(new_n623), .A3(new_n648), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n705), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n653), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n685), .A2(new_n623), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n672), .B(new_n760), .C1(new_n675), .C2(new_n676), .ZN(new_n761));
  NAND2_X1  g560(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n762), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n689), .A2(new_n672), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n652), .A2(new_n552), .A3(new_n647), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n759), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  NAND4_X1  g571(.A1(new_n679), .A2(new_n342), .A3(new_n680), .A4(new_n757), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n342), .A2(new_n553), .A3(new_n647), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n774), .B(new_n778), .C1(new_n770), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n758), .B2(new_n662), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n397), .A2(new_n648), .A3(G99gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT111), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n770), .B2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n515), .A2(new_n648), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n515), .A2(new_n791), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n679), .A2(new_n680), .A3(new_n757), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n785), .A2(new_n786), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n788), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(G106gat), .B1(new_n769), .B2(new_n789), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n795), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(new_n787), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n797), .A2(new_n800), .ZN(G1339gat));
  NAND3_X1  g600(.A1(new_n612), .A2(new_n635), .A3(new_n613), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n629), .B(new_n802), .C1(new_n638), .C2(KEYINPUT10), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n637), .A3(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n630), .C1(new_n633), .C2(new_n636), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT113), .A3(new_n644), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT113), .B1(new_n806), .B2(new_n644), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT55), .B(new_n804), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n646), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n803), .A2(new_n637), .A3(KEYINPUT54), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n644), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n813), .B1(new_n816), .B2(new_n807), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(KEYINPUT114), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n684), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT103), .B1(new_n271), .B2(new_n276), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n811), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n272), .A2(new_n273), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n252), .A3(new_n269), .A4(new_n266), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n203), .B1(new_n268), .B2(new_n262), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n264), .A2(new_n265), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n251), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n827), .A2(new_n647), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n672), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n827), .A2(new_n830), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n822), .A2(new_n834), .A3(new_n811), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n625), .A2(new_n538), .A3(new_n580), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n538), .B1(new_n625), .B2(new_n580), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n730), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n649), .A2(new_n685), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n450), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n653), .A2(new_n342), .A3(new_n397), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n278), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n842), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n847), .A2(new_n451), .A3(new_n735), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n343), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n685), .A2(new_n355), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  NAND4_X1  g650(.A1(new_n848), .A2(new_n349), .A3(new_n343), .A4(new_n647), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n845), .B2(new_n648), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1341gat));
  NOR3_X1   g655(.A1(new_n845), .A2(new_n352), .A3(new_n730), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n849), .A2(new_n730), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n858), .B2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n849), .B2(new_n730), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(G1342gat));
  NAND2_X1  g661(.A1(new_n672), .A2(new_n343), .ZN(new_n863));
  AOI211_X1 g662(.A(G134gat), .B(new_n863), .C1(KEYINPUT117), .C2(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n865), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(KEYINPUT117), .B2(KEYINPUT56), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n843), .A2(new_n672), .A3(new_n844), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(G134gat), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n869), .A2(new_n868), .A3(G134gat), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n866), .B(new_n867), .C1(new_n870), .C2(new_n871), .ZN(G1343gat));
  NAND3_X1  g671(.A1(new_n652), .A2(new_n343), .A3(new_n662), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT119), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n847), .B2(new_n450), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n515), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n819), .A2(new_n820), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n646), .A3(new_n810), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n276), .B2(new_n271), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n582), .B(new_n626), .C1(new_n881), .C2(new_n831), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n623), .B1(new_n882), .B2(new_n838), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(new_n841), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT121), .B(new_n878), .C1(new_n883), .C2(new_n841), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n874), .B1(new_n876), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n278), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n502), .A2(new_n515), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n847), .A2(new_n343), .A3(new_n735), .A4(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(G141gat), .A3(new_n278), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n685), .B(new_n874), .C1(new_n876), .C2(new_n888), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n893), .B1(new_n897), .B2(G141gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(new_n892), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n408), .A3(new_n647), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n647), .B(new_n874), .C1(new_n876), .C2(new_n888), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n902), .A2(new_n903), .A3(G148gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n836), .A2(new_n837), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n822), .A2(new_n811), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n683), .B2(new_n684), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n831), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n623), .B1(new_n908), .B2(new_n838), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n450), .B(new_n875), .C1(new_n909), .C2(new_n841), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n649), .A2(new_n277), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n450), .B1(new_n883), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n877), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n648), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n874), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n901), .B1(new_n904), .B2(new_n916), .ZN(G1345gat));
  INV_X1    g716(.A(new_n416), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n889), .B2(new_n730), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n416), .A3(new_n623), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n889), .B2(new_n905), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n863), .A2(G162gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n847), .A2(new_n735), .A3(new_n891), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n652), .B1(new_n840), .B2(new_n842), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(new_n342), .A3(new_n451), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n685), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n342), .A2(new_n733), .A3(new_n734), .A4(new_n743), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n843), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n278), .A2(new_n285), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  INV_X1    g731(.A(new_n930), .ZN(new_n933));
  OAI21_X1  g732(.A(G176gat), .B1(new_n933), .B2(new_n648), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n927), .A2(new_n286), .A3(new_n647), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND2_X1  g735(.A1(new_n930), .A2(new_n623), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G183gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n289), .A3(new_n623), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n938), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n938), .A2(new_n939), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n941), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n290), .A3(new_n672), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n672), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT61), .B(new_n290), .C1(new_n930), .C2(new_n672), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR3_X1   g750(.A1(new_n502), .A2(new_n343), .A3(new_n515), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n926), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n685), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n733), .A2(new_n342), .A3(new_n662), .A4(new_n734), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n910), .B2(new_n913), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n277), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  INV_X1    g757(.A(G204gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n953), .A2(new_n959), .A3(new_n647), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g761(.A(new_n955), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n914), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n961), .B(new_n962), .C1(new_n959), .C2(new_n964), .ZN(G1353gat));
  INV_X1    g764(.A(G211gat), .ZN(new_n966));
  AOI211_X1 g765(.A(new_n730), .B(new_n955), .C1(new_n910), .C2(new_n913), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(KEYINPUT125), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n956), .A2(new_n623), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n969), .A2(new_n970), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n910), .A2(new_n913), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n977), .A2(KEYINPUT125), .A3(new_n623), .A4(new_n963), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT125), .B1(new_n956), .B2(new_n623), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n975), .B(new_n976), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n926), .A2(new_n966), .A3(new_n623), .A4(new_n952), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n974), .A2(new_n981), .A3(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n953), .B2(new_n672), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n672), .A2(new_n317), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n956), .B2(new_n986), .ZN(G1355gat));
endmodule


