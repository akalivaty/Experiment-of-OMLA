//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT70), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n193), .B(new_n198), .C1(new_n194), .C2(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT66), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G137), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT11), .B1(new_n203), .B2(G134), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n204), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n205), .B2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n202), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n204), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n201), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n200), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT68), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n222), .A2(new_n224), .A3(G116), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n221), .B2(G116), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n220), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n220), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(new_n224), .A3(G116), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n229), .A4(new_n226), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n238), .A2(new_n191), .B1(new_n189), .B2(G128), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n194), .B2(new_n238), .ZN(new_n242));
  AND4_X1   g056(.A1(new_n241), .A2(new_n238), .A3(new_n189), .A4(new_n191), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n206), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n205), .A2(G137), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n219), .A2(new_n236), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n251), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n236), .B1(new_n219), .B2(new_n250), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT28), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT29), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n187), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n246), .A2(new_n249), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n238), .A2(new_n189), .A3(new_n191), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n194), .A2(new_n241), .A3(new_n238), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n239), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n196), .B1(new_n213), .B2(new_n217), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n235), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n253), .B1(new_n251), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n255), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .A4(new_n267), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n219), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n275), .B2(new_n276), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(new_n235), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n251), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n287), .B2(new_n266), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n269), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n251), .A3(new_n267), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n286), .A2(new_n293), .A3(new_n251), .A4(new_n267), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n254), .A2(new_n278), .A3(new_n255), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(new_n267), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(G234), .B2(new_n187), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT16), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n306), .B2(G125), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(G125), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G146), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n317), .A3(new_n188), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n221), .A2(new_n237), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT68), .B(G119), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT23), .B(new_n322), .C1(new_n323), .C2(new_n237), .ZN(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n323), .B2(G128), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n329), .B(new_n322), .C1(new_n323), .C2(new_n237), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n321), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n307), .A2(new_n310), .B1(G125), .B2(new_n306), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n188), .B(new_n314), .C1(new_n336), .C2(new_n305), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n316), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n324), .A2(new_n327), .ZN(new_n339));
  INV_X1    g153(.A(new_n329), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n322), .B1(new_n323), .B2(new_n237), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n339), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT76), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n335), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n316), .A2(new_n320), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n328), .A2(new_n333), .A3(new_n330), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n333), .B1(new_n328), .B2(new_n330), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n338), .A2(new_n342), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n348), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n187), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n349), .B1(new_n335), .B2(new_n343), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n355), .A3(new_n348), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n304), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n303), .A2(G902), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n301), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n370), .A2(KEYINPUT3), .A3(G104), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n370), .B2(G104), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT77), .B1(new_n370), .B2(G104), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n376), .B2(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n370), .A2(KEYINPUT3), .A3(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n374), .A4(new_n377), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(G101), .C1(new_n373), .C2(new_n378), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n200), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n370), .A2(G104), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n376), .A2(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT10), .A3(new_n244), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n385), .A2(new_n392), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(new_n274), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT78), .B(new_n396), .C1(new_n397), .C2(new_n274), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n218), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n395), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n395), .B2(new_n402), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n344), .A2(G227), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n393), .A2(new_n244), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n397), .A2(new_n274), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n218), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n244), .A2(new_n392), .A3(new_n385), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n397), .A2(new_n274), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n395), .A2(new_n402), .A3(new_n403), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n410), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n369), .B1(new_n409), .B2(new_n422), .ZN(new_n423));
  AOI221_X4 g237(.A(new_n414), .B1(new_n213), .B2(new_n217), .C1(new_n416), .C2(new_n417), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT12), .B1(new_n418), .B2(new_n218), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n408), .B1(new_n404), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT78), .B1(new_n416), .B2(new_n396), .ZN(new_n428));
  INV_X1    g242(.A(new_n401), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n389), .A2(new_n394), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n218), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n421), .A3(new_n410), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n433), .A3(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n423), .A2(G469), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n187), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n408), .B1(new_n404), .B2(new_n405), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n420), .A2(new_n421), .A3(new_n410), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n440), .B2(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n344), .A2(G952), .ZN(new_n443));
  NAND2_X1  g257(.A1(G234), .A2(G237), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(G898), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(G902), .A3(G953), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n386), .A2(new_n235), .A3(new_n388), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n233), .A2(KEYINPUT5), .A3(new_n229), .A4(new_n226), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n323), .A2(new_n457), .A3(G116), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(G113), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n393), .A2(new_n234), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G122), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(KEYINPUT6), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n467), .A3(new_n463), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n193), .B(G125), .C1(new_n194), .C2(new_n195), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n274), .B2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n344), .A2(G224), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n462), .B(KEYINPUT8), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(new_n234), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n397), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n477), .B2(new_n460), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n470), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n470), .B2(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n465), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n187), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n454), .B1(new_n473), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n490), .B2(new_n465), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n453), .A3(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n450), .B(new_n452), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n442), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  XNOR2_X1  g312(.A(G113), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n376), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n320), .B1(new_n188), .B2(new_n336), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n502));
  AOI21_X1  g316(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n502), .B2(new_n503), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(KEYINPUT18), .A3(G131), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT82), .B1(new_n509), .B2(new_n245), .ZN(new_n510));
  OR3_X1    g324(.A1(new_n509), .A2(new_n245), .A3(KEYINPUT82), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n501), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT83), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(G131), .C1(new_n502), .C2(new_n503), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n504), .A2(new_n245), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n308), .B1(new_n309), .B2(G140), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n306), .A2(KEYINPUT73), .A3(G125), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n312), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n188), .B1(new_n526), .B2(new_n314), .ZN(new_n527));
  INV_X1    g341(.A(new_n337), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT84), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n316), .A2(new_n530), .A3(new_n337), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n500), .B(new_n513), .C1(new_n522), .C2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT19), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n312), .A2(new_n317), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n336), .B2(new_n534), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n521), .B(new_n316), .C1(G146), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n500), .B1(new_n537), .B2(new_n513), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n498), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  AOI211_X1 g357(.A(KEYINPUT20), .B(new_n543), .C1(new_n533), .C2(new_n539), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n513), .B1(new_n522), .B2(new_n532), .ZN(new_n545));
  INV_X1    g359(.A(new_n500), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n547), .B2(new_n533), .ZN(new_n548));
  INV_X1    g362(.A(G475), .ZN(new_n549));
  OAI22_X1  g363(.A1(new_n542), .A2(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT85), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n513), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n316), .A2(new_n530), .A3(new_n337), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n530), .B1(new_n316), .B2(new_n337), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n521), .A2(new_n519), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n515), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n538), .B1(new_n560), .B2(new_n500), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT20), .B1(new_n561), .B2(new_n543), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n540), .A2(new_n498), .A3(new_n541), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n533), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n556), .A2(new_n559), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n500), .B1(new_n566), .B2(new_n513), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n187), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G475), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n569), .A3(KEYINPUT85), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n190), .A2(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n237), .A2(G143), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n205), .ZN(new_n574));
  XNOR2_X1  g388(.A(G116), .B(G122), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n370), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n228), .A2(KEYINPUT14), .A3(G122), .ZN(new_n577));
  INV_X1    g391(.A(new_n575), .ZN(new_n578));
  OAI211_X1 g392(.A(G107), .B(new_n577), .C1(new_n578), .C2(KEYINPUT14), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n571), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n581), .A2(KEYINPUT13), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n572), .B1(new_n581), .B2(KEYINPUT13), .ZN(new_n583));
  OAI21_X1  g397(.A(G134), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n573), .A2(new_n205), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n575), .B(new_n370), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n495), .A2(new_n302), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n187), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n593), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n552), .A2(new_n570), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n368), .A2(new_n497), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT88), .B(G101), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G3));
  NAND2_X1  g415(.A1(new_n292), .A2(new_n294), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n267), .B1(new_n256), .B2(new_n279), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n187), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n604), .A2(G472), .B1(new_n296), .B2(new_n298), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n442), .A2(new_n605), .A3(new_n367), .A4(new_n496), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n489), .A2(new_n493), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(new_n451), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT89), .B(new_n452), .C1(new_n489), .C2(new_n493), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n449), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n552), .A2(new_n570), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n588), .A2(new_n590), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(KEYINPUT90), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n591), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n591), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(G478), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n594), .A2(new_n187), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n619), .B(new_n621), .C1(G478), .C2(new_n592), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT91), .B1(new_n613), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n625), .B(new_n622), .C1(new_n552), .C2(new_n570), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n612), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT92), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n612), .B(KEYINPUT92), .C1(new_n624), .C2(new_n626), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n606), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT94), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n548), .A2(new_n634), .A3(new_n549), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT94), .B1(new_n568), .B2(G475), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n542), .B2(new_n544), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT93), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n593), .B(new_n595), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n606), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT96), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n354), .A2(new_n355), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n365), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n651), .B1(new_n364), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n604), .A2(G472), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT25), .B1(new_n362), .B2(new_n187), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n358), .B(G902), .C1(new_n360), .C2(new_n361), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n303), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n365), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(KEYINPUT97), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n296), .A2(new_n298), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n656), .A2(new_n657), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n497), .A2(new_n664), .A3(new_n598), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n442), .A2(new_n496), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n445), .B(KEYINPUT98), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(G900), .B2(new_n448), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n637), .A2(new_n641), .A3(new_n642), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n491), .A2(new_n453), .A3(new_n492), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n453), .B1(new_n491), .B2(new_n492), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n451), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT89), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n608), .A2(new_n607), .A3(new_n451), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G472), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n259), .A2(new_n280), .A3(new_n281), .ZN(new_n680));
  INV_X1    g494(.A(new_n268), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n282), .A2(new_n288), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n663), .A2(KEYINPUT32), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n656), .A2(new_n662), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n672), .A2(new_n678), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  AOI21_X1  g505(.A(new_n597), .B1(new_n552), .B2(new_n570), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n608), .B(new_n694), .ZN(new_n695));
  OR3_X1    g509(.A1(new_n693), .A2(new_n695), .A3(new_n452), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n364), .A2(new_n655), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n685), .A2(new_n686), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n287), .A2(new_n267), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n257), .A2(new_n258), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n699), .B(new_n187), .C1(new_n267), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G472), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT100), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  INV_X1    g518(.A(new_n702), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n704), .B(new_n705), .C1(new_n685), .C2(new_n686), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n697), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n496), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n435), .B2(new_n441), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n670), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n696), .A2(new_n707), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n190), .ZN(G45));
  INV_X1    g530(.A(new_n670), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n622), .B(new_n717), .C1(new_n552), .C2(new_n570), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n689), .A2(new_n718), .A3(new_n709), .A4(new_n678), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  AOI21_X1  g534(.A(new_n410), .B1(new_n432), .B2(new_n421), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n420), .A2(new_n421), .A3(new_n410), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n187), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n436), .B(new_n187), .C1(new_n721), .C2(new_n722), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(KEYINPUT102), .A3(new_n725), .ZN(new_n726));
  OR3_X1    g540(.A1(new_n440), .A2(KEYINPUT102), .A3(new_n436), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n301), .A2(new_n728), .A3(new_n367), .A4(new_n496), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n629), .B2(new_n630), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT41), .B(G113), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n644), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NOR3_X1   g549(.A1(new_n364), .A2(new_n651), .A3(new_n655), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT97), .B1(new_n660), .B2(new_n661), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n678), .A2(new_n738), .A3(new_n301), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n552), .A2(new_n570), .A3(new_n597), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n450), .B(new_n708), .C1(new_n726), .C2(new_n727), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(KEYINPUT103), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n708), .B1(new_n726), .B2(new_n727), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n740), .A3(new_n449), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n678), .A2(new_n738), .A3(new_n301), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  NAND3_X1  g563(.A1(new_n728), .A2(new_n449), .A3(new_n496), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n292), .B(new_n294), .C1(new_n680), .C2(new_n267), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n298), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n679), .B1(new_n296), .B2(new_n187), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n367), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n692), .A2(new_n678), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NOR3_X1   g574(.A1(new_n753), .A2(new_n697), .A3(new_n754), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n718), .A2(new_n678), .A3(new_n744), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(new_n368), .ZN(new_n764));
  AOI211_X1 g578(.A(G469), .B(G902), .C1(new_n438), .C2(new_n439), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n427), .A2(new_n433), .A3(G469), .ZN(new_n766));
  INV_X1    g580(.A(new_n437), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n496), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT104), .B(new_n496), .C1(new_n765), .C2(new_n768), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n489), .A2(new_n451), .A3(new_n493), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(KEYINPUT105), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n773), .B1(new_n769), .B2(new_n770), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT105), .B1(new_n776), .B2(new_n772), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n764), .B(new_n718), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n431), .B1(new_n400), .B2(new_n401), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n408), .B1(new_n783), .B2(new_n403), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n420), .A2(new_n421), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n432), .A2(new_n784), .B1(new_n785), .B2(new_n408), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n437), .B1(new_n786), .B2(G469), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n708), .B1(new_n787), .B2(new_n725), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n774), .B1(new_n788), .B2(KEYINPUT104), .ZN(new_n789));
  INV_X1    g603(.A(new_n772), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n782), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n776), .A2(KEYINPUT105), .A3(new_n772), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(KEYINPUT106), .A3(new_n764), .A4(new_n718), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n780), .A2(new_n781), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n613), .A2(new_n623), .A3(new_n670), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n368), .B(new_n796), .C1(new_n791), .C2(new_n792), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT107), .B1(new_n797), .B2(KEYINPUT42), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n780), .A2(KEYINPUT107), .A3(new_n794), .A4(new_n781), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n671), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n793), .A2(new_n764), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NOR2_X1   g620(.A1(new_n550), .A2(new_n551), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT85), .B1(new_n564), .B2(new_n569), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n623), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT110), .B1(new_n810), .B2(KEYINPUT109), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT43), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n810), .B2(KEYINPUT110), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n605), .ZN(new_n816));
  INV_X1    g630(.A(new_n697), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT45), .B1(new_n423), .B2(new_n434), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n436), .B(new_n822), .C1(KEYINPUT45), .C2(new_n786), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT46), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n823), .A2(new_n824), .A3(new_n437), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n823), .B2(new_n437), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n725), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(new_n496), .A3(new_n711), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n774), .A3(new_n821), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G137), .ZN(G39));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n496), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT47), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(KEYINPUT47), .A3(new_n496), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n796), .A2(new_n301), .A3(new_n367), .A4(new_n773), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT111), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  NAND3_X1  g653(.A1(new_n367), .A2(new_n451), .A3(new_n496), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n809), .B(new_n623), .C1(KEYINPUT112), .C2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(KEYINPUT112), .B2(new_n840), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT113), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n702), .B1(new_n299), .B2(new_n300), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n704), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n698), .A2(KEYINPUT100), .A3(new_n702), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n728), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n695), .B1(new_n728), .B2(new_n849), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n850), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n843), .A2(new_n848), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n757), .A2(new_n758), .B1(new_n729), .B2(new_n644), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n494), .B(new_n623), .C1(new_n807), .C2(new_n808), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n606), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n599), .A2(new_n665), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n552), .A2(new_n570), .A3(new_n642), .ZN(new_n861));
  INV_X1    g675(.A(new_n494), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT115), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n645), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n748), .A2(new_n857), .A3(new_n860), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n731), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n817), .A2(new_n657), .A3(new_n752), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n796), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n793), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n637), .A2(new_n641), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n642), .A2(new_n773), .A3(new_n717), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n689), .A2(new_n709), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n805), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n799), .A2(new_n867), .A3(new_n800), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n690), .A2(new_n719), .A3(new_n762), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n670), .B(KEYINPUT116), .Z(new_n879));
  AND2_X1   g693(.A1(new_n788), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n678), .A3(new_n692), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n707), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT52), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n744), .A2(new_n678), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n884), .A2(new_n869), .B1(new_n739), .B2(new_n672), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n847), .A2(new_n758), .A3(new_n697), .A4(new_n880), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n719), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n690), .A2(new_n762), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n883), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n866), .A2(new_n874), .A3(new_n731), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n799), .A3(new_n891), .A4(new_n800), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT119), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n883), .A2(new_n888), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n883), .B2(new_n888), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n801), .A3(new_n893), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n799), .A2(new_n867), .A3(new_n800), .A4(new_n875), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n883), .A2(new_n888), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n901), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n899), .B(new_n895), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n897), .B(new_n898), .C1(new_n906), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n894), .A2(new_n895), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n905), .B2(new_n895), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n913), .B2(new_n917), .ZN(new_n919));
  INV_X1    g733(.A(new_n669), .ZN(new_n920));
  INV_X1    g734(.A(new_n756), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n815), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n496), .B1(new_n726), .B2(new_n727), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n774), .B(new_n923), .C1(new_n835), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n744), .A2(new_n452), .A3(new_n695), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT121), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(KEYINPUT50), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT50), .ZN(new_n929));
  INV_X1    g743(.A(new_n927), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n744), .A2(new_n774), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n815), .A2(new_n920), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n445), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n848), .A2(new_n367), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n809), .A2(new_n622), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n936), .A2(KEYINPUT122), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT122), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n934), .A2(new_n761), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n925), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT51), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n624), .A2(new_n626), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n884), .ZN(new_n946));
  OAI221_X1 g760(.A(new_n443), .B1(new_n945), .B2(new_n936), .C1(new_n922), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n934), .A2(new_n764), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n941), .A2(KEYINPUT123), .A3(new_n942), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT123), .B1(new_n941), .B2(new_n942), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n943), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n918), .A2(new_n919), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(G952), .A2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n856), .B1(new_n956), .B2(new_n957), .ZN(G75));
  NAND2_X1  g772(.A1(new_n466), .A2(new_n468), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n472), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n895), .B1(new_n907), .B2(new_n910), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT118), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n963), .A2(new_n911), .B1(new_n892), .B2(new_n896), .ZN(new_n964));
  INV_X1    g778(.A(G210), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n187), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(KEYINPUT56), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n344), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n966), .A2(KEYINPUT56), .A3(new_n961), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G51));
  XNOR2_X1  g786(.A(new_n437), .B(KEYINPUT124), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT57), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n963), .A2(new_n911), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n975), .A2(new_n898), .A3(new_n897), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n898), .B1(new_n975), .B2(new_n897), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n721), .B2(new_n722), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n964), .A2(new_n187), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n823), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n968), .B1(new_n979), .B2(new_n981), .ZN(G54));
  AND2_X1   g796(.A1(KEYINPUT58), .A2(G475), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n980), .A2(new_n540), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n540), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(new_n968), .ZN(G60));
  AND2_X1   g800(.A1(new_n617), .A2(new_n618), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n620), .B(KEYINPUT59), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n976), .B2(new_n977), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n969), .ZN(new_n991));
  INV_X1    g805(.A(new_n988), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n918), .B2(new_n919), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(new_n987), .ZN(G63));
  XNOR2_X1  g808(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n302), .A2(new_n187), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n964), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n654), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n361), .B(new_n360), .C1(new_n964), .C2(new_n998), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n969), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT61), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1000), .A2(KEYINPUT61), .A3(new_n969), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G66));
  NAND2_X1  g820(.A1(new_n447), .A2(G224), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n867), .B2(G953), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n959), .B1(G898), .B2(new_n344), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(G69));
  NAND2_X1  g826(.A1(new_n283), .A2(new_n285), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(new_n536), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(G900), .B2(G953), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n828), .A2(new_n764), .A3(new_n758), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n719), .A2(new_n1018), .A3(new_n805), .A4(new_n885), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n838), .A2(new_n829), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n801), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1017), .B1(new_n1022), .B2(new_n344), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n344), .B1(G227), .B2(G900), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n715), .A2(new_n878), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT62), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n712), .A2(new_n773), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n861), .B1(new_n809), .B2(new_n622), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n764), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n838), .A2(new_n829), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n344), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n1015), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1024), .A2(new_n1026), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1036), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1025), .B1(new_n1038), .B2(new_n1023), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1037), .A2(new_n1039), .ZN(G72));
  NOR2_X1   g854(.A1(new_n287), .A2(new_n267), .ZN(new_n1041));
  NOR4_X1   g855(.A1(new_n1020), .A2(new_n731), .A3(new_n1021), .A4(new_n866), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n699), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1047), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n916), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(KEYINPUT127), .ZN(new_n1050));
  INV_X1    g864(.A(new_n867), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1044), .B1(new_n1034), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n968), .B1(new_n1052), .B2(new_n1047), .ZN(new_n1053));
  AND3_X1   g867(.A1(new_n1046), .A2(new_n1050), .A3(new_n1053), .ZN(G57));
endmodule


