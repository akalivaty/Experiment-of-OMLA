//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  XOR2_X1   g000(.A(KEYINPUT87), .B(G475), .Z(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(new_n188), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT74), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n188), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G237), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G214), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(G237), .A2(G953), .ZN(new_n202));
  AOI21_X1  g016(.A(G143), .B1(new_n202), .B2(G214), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT18), .B(G131), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(new_n200), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT18), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n196), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G113), .B(G122), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(KEYINPUT85), .ZN(new_n215));
  INV_X1    g029(.A(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  INV_X1    g031(.A(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G146), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(G146), .B1(new_n220), .B2(new_n221), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n201), .B2(new_n203), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n208), .A3(new_n206), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n226), .A2(KEYINPUT86), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT17), .B(G131), .C1(new_n201), .C2(new_n203), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n211), .B(new_n215), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n211), .B1(new_n231), .B2(new_n234), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n214), .B1(new_n237), .B2(KEYINPUT88), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n211), .B(new_n239), .C1(new_n234), .C2(new_n231), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n187), .B1(new_n241), .B2(G902), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT19), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n188), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n222), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n226), .A2(new_n228), .ZN(new_n250));
  OAI22_X1  g064(.A1(new_n249), .A2(new_n250), .B1(new_n196), .B2(new_n210), .ZN(new_n251));
  INV_X1    g065(.A(new_n214), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n235), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT20), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n258), .A3(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n242), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G952), .ZN(new_n262));
  AOI211_X1 g076(.A(G953), .B(new_n262), .C1(G234), .C2(G237), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  AOI211_X1 g078(.A(new_n264), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT21), .B(G898), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n200), .A2(G128), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT13), .Z(new_n269));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n200), .B2(G128), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT89), .A3(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(G134), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n277), .A3(new_n268), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT78), .B(G107), .ZN(new_n279));
  XNOR2_X1  g093(.A(G116), .B(G122), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n276), .B(new_n278), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n284));
  INV_X1    g098(.A(new_n278), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n274), .B2(new_n268), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n268), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G134), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT90), .A3(new_n278), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT14), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G107), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G122), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n295), .B2(KEYINPUT14), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n282), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n283), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  INV_X1    g114(.A(G217), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(G953), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n283), .A2(new_n298), .A3(new_n302), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n307));
  INV_X1    g121(.A(G478), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT15), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n283), .A2(new_n298), .A3(new_n302), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n302), .B1(new_n283), .B2(new_n298), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n307), .B(new_n264), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n261), .A2(new_n267), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n294), .A2(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT2), .B(G113), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n293), .A2(G104), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n279), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n293), .A2(G104), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT79), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n335), .A2(G101), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n327), .A2(new_n333), .A3(new_n336), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n336), .B1(new_n327), .B2(new_n333), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(new_n333), .A3(new_n342), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT4), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n324), .B(new_n339), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n331), .B1(new_n279), .B2(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G101), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n350));
  INV_X1    g164(.A(G113), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT5), .ZN(new_n353));
  INV_X1    g167(.A(new_n322), .ZN(new_n354));
  INV_X1    g168(.A(new_n323), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n346), .A2(new_n359), .A3(new_n357), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n245), .A2(new_n247), .A3(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n200), .A2(KEYINPUT65), .A3(G146), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT65), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n189), .B2(G143), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n272), .B1(new_n364), .B2(KEYINPUT1), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n200), .A2(G146), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n248), .B2(new_n200), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n218), .B(new_n369), .C1(new_n370), .C2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n371), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n191), .B2(G143), .ZN(new_n376));
  AND2_X1   g190(.A1(KEYINPUT0), .A2(G128), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n377), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n218), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n198), .A2(G224), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n358), .A2(new_n386), .A3(new_n360), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n363), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n344), .A2(new_n348), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n356), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n359), .B(KEYINPUT8), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n353), .A2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n352), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n354), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n394), .A2(new_n395), .B1(new_n354), .B2(new_n355), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n390), .B(new_n391), .C1(new_n396), .C2(new_n389), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  INV_X1    g212(.A(new_n382), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n384), .A4(new_n373), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n374), .B2(new_n382), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n398), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n362), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(new_n400), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT84), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n388), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n388), .B2(new_n407), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n317), .B(new_n318), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G221), .ZN(new_n415));
  INV_X1    g229(.A(new_n300), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(new_n264), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n419));
  OAI21_X1  g233(.A(G128), .B1(new_n371), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n245), .A2(new_n247), .A3(G143), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n367), .A2(new_n365), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT81), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n369), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n349), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n389), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n380), .A2(new_n381), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(new_n339), .C1(new_n343), .C2(new_n345), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT68), .A2(G131), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n277), .A2(G137), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT11), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT66), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT11), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G137), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G134), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n439), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT11), .A2(G134), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT67), .B1(new_n448), .B2(G137), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n445), .A3(KEYINPUT11), .A4(G134), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n437), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n441), .A2(new_n443), .B1(new_n277), .B2(G137), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n437), .C1(new_n454), .C2(new_n438), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n436), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n428), .A2(new_n429), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n430), .A2(new_n431), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n435), .A2(new_n460), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n198), .A2(G227), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n421), .A2(new_n422), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n423), .A2(new_n424), .B1(new_n468), .B2(new_n368), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n389), .B1(new_n469), .B2(new_n426), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n431), .B1(new_n344), .B2(new_n348), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n431), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n389), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n428), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT12), .A3(new_n458), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n466), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n462), .A3(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(G469), .B(G902), .C1(new_n467), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G469), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT12), .B1(new_n477), .B2(new_n458), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n473), .B(new_n457), .C1(new_n428), .C2(new_n476), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n462), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n466), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n459), .A2(new_n462), .A3(new_n480), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n489), .B2(new_n264), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n418), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n414), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n452), .B(new_n208), .C1(new_n454), .C2(new_n438), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n438), .B2(new_n446), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n475), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n434), .B1(new_n456), .B2(new_n453), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n431), .A2(KEYINPUT69), .A3(new_n495), .A4(new_n494), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n495), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n431), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n498), .A3(KEYINPUT30), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n324), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n202), .A2(G210), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT27), .Z(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G101), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n324), .B(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n498), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n508), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT31), .ZN(new_n517));
  INV_X1    g331(.A(new_n512), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT28), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n500), .A2(new_n324), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n519), .B1(new_n525), .B2(new_n515), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n518), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT31), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n508), .A2(new_n528), .A3(new_n512), .A4(new_n515), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n512), .B1(new_n524), .B2(new_n526), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n508), .A2(new_n518), .A3(new_n515), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n515), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT72), .B1(new_n515), .B2(new_n519), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT73), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n542), .A3(new_n523), .ZN(new_n543));
  INV_X1    g357(.A(new_n515), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n514), .B1(new_n506), .B2(new_n498), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT28), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n512), .A2(KEYINPUT29), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n543), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n538), .A2(new_n549), .A3(G902), .ZN(new_n550));
  INV_X1    g364(.A(G472), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n534), .B(new_n535), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n301), .B1(G234), .B2(new_n264), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n193), .A2(new_n195), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n319), .B2(G128), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n272), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(new_n561), .C1(G119), .C2(new_n272), .ZN(new_n562));
  XNOR2_X1  g376(.A(G119), .B(G128), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT24), .B(G110), .Z(new_n564));
  OAI22_X1  g378(.A1(new_n562), .A2(G110), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n222), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n562), .A2(G110), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n223), .B2(new_n224), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n572), .A3(new_n568), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n571), .A2(new_n577), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n557), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n555), .A2(new_n556), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n554), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI221_X1 g397(.A(new_n557), .B1(new_n555), .B2(new_n556), .C1(new_n579), .C2(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n553), .A2(G902), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n579), .B2(new_n580), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n492), .A2(new_n552), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT92), .B(G101), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G3));
  NAND2_X1  g406(.A1(new_n530), .A2(new_n264), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n532), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n595), .A2(new_n588), .A3(new_n491), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n388), .A2(new_n407), .A3(new_n408), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n408), .B1(new_n388), .B2(new_n407), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n318), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G478), .A2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n306), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(G478), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n312), .A2(new_n313), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT33), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(G478), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n261), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n599), .A2(new_n267), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND3_X1  g424(.A1(new_n242), .A2(new_n316), .A3(new_n260), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n599), .A2(new_n267), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n596), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(new_n595), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n569), .B(new_n617), .Z(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n586), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n585), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n621), .B(new_n418), .C1(new_n482), .C2(new_n490), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n412), .A2(new_n413), .ZN(new_n624));
  INV_X1    g438(.A(new_n318), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n623), .A3(new_n626), .A4(new_n317), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT93), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n388), .A2(new_n407), .ZN(new_n632));
  INV_X1    g446(.A(new_n408), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n388), .A2(new_n407), .A3(new_n408), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n263), .B1(new_n265), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n316), .A2(new_n242), .A3(new_n260), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n631), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n640), .B(new_n318), .C1(new_n597), .C2(new_n598), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(KEYINPUT94), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n552), .B(new_n623), .C1(new_n641), .C2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  XOR2_X1   g459(.A(new_n638), .B(KEYINPUT39), .Z(new_n646));
  OAI211_X1 g460(.A(new_n418), .B(new_n646), .C1(new_n482), .C2(new_n490), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT96), .Z(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n314), .A2(new_n309), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n318), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n260), .B2(new_n242), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n583), .A2(new_n584), .B1(new_n586), .B2(new_n619), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT95), .Z(new_n657));
  NOR2_X1   g471(.A1(new_n544), .A2(new_n545), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n658), .B2(new_n518), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n518), .B1(new_n508), .B2(new_n515), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n534), .A2(new_n535), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n624), .B(KEYINPUT38), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n657), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n649), .A2(new_n650), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  NAND3_X1  g482(.A1(new_n605), .A2(new_n261), .A3(new_n639), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n599), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n552), .A2(new_n623), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT97), .B(G146), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G48));
  NAND2_X1  g487(.A1(new_n467), .A2(new_n481), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n264), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n483), .A3(new_n264), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n418), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n552), .A2(new_n607), .A3(new_n589), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n552), .A2(new_n612), .A3(new_n589), .A4(new_n678), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  AND2_X1   g497(.A1(new_n636), .A2(new_n317), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n552), .A2(new_n684), .A3(new_n621), .A4(new_n678), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  INV_X1    g500(.A(new_n267), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n676), .A2(new_n418), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n634), .A2(new_n635), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT101), .B1(new_n689), .B2(new_n654), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n654), .B(KEYINPUT101), .C1(new_n597), .C2(new_n598), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n517), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n512), .B1(new_n695), .B2(KEYINPUT98), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n541), .A2(new_n543), .A3(new_n697), .A4(new_n546), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT99), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n529), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI211_X1 g515(.A(KEYINPUT99), .B(new_n694), .C1(new_n696), .C2(new_n698), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n531), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n588), .B(KEYINPUT100), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n693), .A2(new_n594), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND4_X1  g520(.A1(new_n676), .A2(new_n418), .A3(new_n677), .A4(new_n621), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n707), .A2(new_n599), .A3(new_n669), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n703), .A2(new_n594), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NAND2_X1  g524(.A1(new_n535), .A2(KEYINPUT103), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n530), .A2(new_n712), .A3(KEYINPUT32), .A4(new_n531), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n534), .A2(KEYINPUT104), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n536), .A2(new_n537), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n264), .B(new_n548), .C1(new_n716), .C2(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT32), .B1(new_n530), .B2(new_n531), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n714), .A2(new_n715), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n413), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n318), .A3(new_n411), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n491), .A2(new_n724), .A3(new_n669), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n722), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n491), .A2(new_n724), .ZN(new_n727));
  INV_X1    g541(.A(new_n669), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n552), .A2(new_n727), .A3(new_n589), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  AND3_X1   g547(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n719), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n588), .B1(new_n735), .B2(new_n718), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n640), .A3(new_n727), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n605), .A2(new_n260), .A3(new_n242), .ZN(new_n743));
  MUX2_X1   g557(.A(new_n740), .B(new_n742), .S(new_n743), .Z(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n595), .A3(new_n621), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n724), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n483), .A2(new_n264), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n483), .B1(new_n489), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n480), .B1(new_n479), .B2(new_n462), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n462), .A2(new_n480), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n457), .B1(new_n432), .B2(new_n435), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n754), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n753), .A3(new_n756), .A4(G469), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n752), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(G469), .A3(new_n756), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT105), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n751), .B1(new_n769), .B2(new_n763), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n482), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT46), .B(new_n752), .C1(new_n757), .C2(new_n764), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n772), .A3(new_n677), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n418), .B(new_n646), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT107), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n766), .B(new_n751), .C1(new_n769), .C2(new_n763), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT106), .B1(new_n779), .B2(new_n482), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n775), .A3(new_n767), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n418), .A4(new_n646), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n750), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n445), .ZN(G39));
  NOR4_X1   g599(.A1(new_n552), .A2(new_n589), .A3(new_n669), .A4(new_n724), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n774), .A2(new_n677), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(KEYINPUT106), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n787), .B(new_n417), .C1(new_n790), .C2(new_n775), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT47), .B1(new_n781), .B2(new_n418), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n655), .A2(new_n639), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n491), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n692), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n797), .B(new_n663), .C1(new_n798), .C2(new_n690), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n644), .A2(new_n671), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n800), .B2(new_n709), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n622), .B1(new_n735), .B2(new_n718), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n636), .A2(new_n631), .A3(new_n640), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n642), .A2(KEYINPUT94), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n805), .B2(new_n670), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n709), .A2(new_n806), .A3(KEYINPUT112), .A4(new_n799), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n795), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n261), .A2(new_n316), .A3(new_n638), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n724), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n552), .A2(new_n623), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT111), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n802), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n703), .A2(new_n594), .A3(new_n621), .A4(new_n725), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n732), .A2(new_n816), .A3(new_n737), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n491), .A2(new_n588), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n267), .B1(new_n606), .B2(new_n611), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n616), .A2(new_n819), .A3(new_n626), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n627), .A2(new_n821), .A3(new_n590), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n685), .A2(new_n679), .A3(new_n682), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n705), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n644), .A2(new_n671), .A3(new_n799), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n703), .A2(new_n594), .A3(new_n708), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n809), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n827), .B2(new_n828), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n809), .A2(new_n825), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n823), .A2(new_n705), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n705), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n818), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n809), .A2(new_n842), .A3(new_n844), .A4(new_n834), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n824), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n732), .A2(new_n737), .A3(new_n816), .A4(new_n817), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(new_n829), .B2(new_n807), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n833), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n837), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n703), .A2(new_n594), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n704), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n744), .A2(new_n263), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n678), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n599), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n676), .A2(new_n677), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n724), .A3(new_n417), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n722), .A2(new_n704), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n589), .A2(new_n864), .A3(new_n664), .A4(new_n263), .ZN(new_n869));
  INV_X1    g683(.A(new_n606), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n262), .B(G953), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n859), .A2(new_n860), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n791), .A2(new_n792), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n863), .A2(new_n418), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n748), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n858), .A2(new_n621), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n605), .A2(new_n261), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n877), .A2(new_n865), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n665), .A2(new_n625), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n861), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT50), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT50), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n861), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n876), .B(new_n879), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n862), .B(new_n872), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n857), .B(new_n887), .C1(new_n886), .C2(new_n885), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n262), .A2(new_n198), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n665), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n743), .B(new_n891), .C1(KEYINPUT49), .C2(new_n863), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n704), .A2(new_n418), .A3(new_n318), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT109), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n863), .A2(KEYINPUT49), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT110), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n894), .A3(new_n664), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(new_n897), .ZN(G75));
  AND3_X1   g712(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT113), .B1(new_n831), .B2(new_n833), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n845), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(G210), .A3(G902), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n363), .A2(new_n387), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n385), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n902), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n902), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n198), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n751), .B(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n855), .A2(new_n856), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n856), .B(new_n845), .C1(new_n899), .C2(new_n900), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n674), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n901), .A2(G902), .A3(new_n763), .A4(new_n769), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n901), .A2(G902), .A3(new_n254), .A4(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT116), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n901), .A2(G902), .A3(new_n920), .ZN(new_n923));
  INV_X1    g737(.A(new_n254), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n910), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(KEYINPUT116), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n914), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n604), .B(KEYINPUT117), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n600), .B(KEYINPUT59), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n910), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n931), .C1(new_n857), .C2(new_n932), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n914), .B2(new_n836), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT118), .B1(new_n937), .B2(new_n930), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n301), .A2(new_n264), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n901), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n579), .A2(new_n580), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n910), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n618), .B(KEYINPUT120), .Z(new_n947));
  NAND3_X1  g761(.A1(new_n901), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  INV_X1    g767(.A(new_n266), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n198), .B1(new_n954), .B2(G224), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n824), .B2(new_n198), .ZN(new_n956));
  INV_X1    g770(.A(G898), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n903), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  NAND2_X1  g773(.A1(new_n778), .A2(new_n783), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n691), .A2(new_n692), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n866), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT124), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n965), .B(new_n962), .C1(new_n778), .C2(new_n783), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n750), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n960), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n732), .A2(new_n737), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n709), .A2(new_n806), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n969), .A2(new_n793), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n967), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n417), .B1(new_n790), .B2(new_n775), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n782), .B1(new_n977), .B2(new_n646), .ZN(new_n978));
  INV_X1    g792(.A(new_n783), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n963), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n965), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n960), .A2(KEYINPUT124), .A3(new_n963), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n793), .A2(new_n970), .A3(new_n973), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n784), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT125), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n198), .B1(new_n976), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n502), .A2(new_n507), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n244), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n637), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT123), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n973), .A2(new_n667), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n606), .A2(new_n611), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT122), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n647), .A2(new_n724), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n736), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n793), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n973), .A2(new_n667), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n996), .A2(new_n1001), .A3(new_n969), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n198), .A3(new_n990), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n992), .A2(KEYINPUT126), .A3(new_n994), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g822(.A(new_n991), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n975), .B1(new_n967), .B2(new_n974), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n985), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n1012), .B2(new_n198), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1005), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1007), .B(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1006), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n1004), .B2(new_n824), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n661), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1010), .A2(new_n1011), .A3(new_n847), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n537), .B1(new_n1022), .B2(new_n1018), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n832), .A2(new_n835), .ZN(new_n1024));
  INV_X1    g838(.A(new_n661), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n537), .A3(new_n1018), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n946), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1021), .A2(new_n1023), .A3(new_n1027), .ZN(G57));
endmodule


