//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n202), .A3(new_n206), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT74), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n211), .A2(new_n212), .A3(new_n207), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  INV_X1    g014(.A(G120gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G113gat), .ZN(new_n217));
  INV_X1    g016(.A(G113gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G120gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT1), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(G134gat), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(G134gat), .B1(new_n222), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n215), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n220), .B(new_n221), .ZN(new_n227));
  INV_X1    g026(.A(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n222), .A2(G134gat), .A3(new_n223), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT75), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n211), .A2(new_n207), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n226), .A3(new_n231), .A4(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n232), .A3(new_n230), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n237));
  OR2_X1    g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n231), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n210), .A2(new_n213), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n236), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n243), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n224), .A2(new_n225), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n237), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n235), .A2(new_n251), .A3(new_n242), .A4(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(KEYINPUT5), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256));
  XNOR2_X1  g055(.A(G57gat), .B(G85gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n243), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n242), .B(new_n236), .C1(new_n246), .C2(new_n247), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT39), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT39), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n267), .A3(new_n243), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n260), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(KEYINPUT80), .A3(new_n260), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT40), .ZN(new_n275));
  INV_X1    g074(.A(new_n272), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT80), .B1(new_n268), .B2(new_n260), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT40), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT81), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n262), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G64gat), .B(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(G36gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT73), .ZN(new_n284));
  INV_X1    g083(.A(G8gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n288));
  INV_X1    g087(.A(G211gat), .ZN(new_n289));
  INV_X1    g088(.A(G218gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT66), .B(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G183gat), .ZN(new_n301));
  OR3_X1    g100(.A1(new_n301), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT27), .B1(new_n301), .B2(KEYINPUT67), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n299), .A2(new_n300), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n309), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n312), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT65), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n306), .B(KEYINPUT24), .Z(new_n327));
  NOR2_X1   g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n297), .A2(G183gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT25), .B1(new_n331), .B2(new_n327), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n320), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G226gat), .ZN(new_n336));
  INV_X1    g135(.A(G233gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n330), .A2(new_n334), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n340), .B2(new_n320), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n295), .B(new_n339), .C1(new_n341), .C2(new_n338), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n338), .B1(new_n335), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n338), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n340), .B2(new_n320), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n294), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n342), .A2(new_n347), .A3(KEYINPUT72), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT72), .B1(new_n342), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n286), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n286), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(KEYINPUT30), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n273), .A2(KEYINPUT40), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n352), .A2(KEYINPUT30), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n281), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358));
  INV_X1    g157(.A(new_n262), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT6), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n245), .A2(new_n254), .A3(new_n260), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n262), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n361), .B2(new_n262), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n364), .B2(new_n358), .ZN(new_n365));
  INV_X1    g164(.A(new_n342), .ZN(new_n366));
  INV_X1    g165(.A(new_n347), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT37), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n351), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT37), .B1(new_n348), .B2(new_n349), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n372), .A2(KEYINPUT38), .B1(new_n351), .B2(new_n368), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT38), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n370), .B(new_n374), .C1(new_n369), .C2(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n365), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n353), .A2(new_n355), .A3(new_n354), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n274), .B1(new_n273), .B2(KEYINPUT40), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n278), .A2(KEYINPUT81), .A3(new_n279), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n359), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G228gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n232), .B2(new_n233), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n294), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n233), .B1(new_n294), .B2(KEYINPUT29), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n213), .B2(new_n210), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n386), .B(new_n337), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n387), .A2(new_n295), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n294), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n293), .B1(new_n291), .B2(new_n287), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n397), .B2(KEYINPUT78), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI221_X1 g198(.A(new_n394), .B1(new_n386), .B2(new_n337), .C1(new_n232), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT31), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n390), .A2(new_n392), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(G228gat), .A3(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT31), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n406));
  XOR2_X1   g205(.A(G78gat), .B(G106gat), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n402), .B2(new_n406), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n385), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n402), .A2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n407), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n384), .A3(new_n409), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n335), .B1(new_n224), .B2(new_n225), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n340), .A2(new_n250), .A3(new_n320), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G227gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(new_n337), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT69), .B(G71gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G99gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(KEYINPUT70), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT33), .B1(new_n427), .B2(KEYINPUT70), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n420), .A2(new_n422), .B1(new_n417), .B2(KEYINPUT33), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(new_n427), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n418), .B(new_n419), .C1(new_n421), .C2(new_n337), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n435), .A2(KEYINPUT71), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n435), .B2(KEYINPUT71), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n431), .A2(new_n433), .B1(new_n438), .B2(new_n437), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT36), .B1(new_n440), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n383), .A2(new_n416), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n353), .A2(new_n355), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n365), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n440), .A2(KEYINPUT84), .A3(new_n441), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT84), .B1(new_n440), .B2(new_n441), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n416), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n442), .A2(new_n416), .A3(new_n443), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(new_n441), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n416), .A2(KEYINPUT35), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n447), .B(new_n364), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n459));
  INV_X1    g258(.A(G29gat), .ZN(new_n460));
  INV_X1    g259(.A(G36gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G50gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G43gat), .ZN(new_n470));
  INV_X1    g269(.A(G43gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G50gat), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT15), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n471), .A2(G50gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n469), .A2(G43gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT15), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n467), .A4(new_n464), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(G1gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT16), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n285), .C1(G1gat), .C2(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(G15gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(G22gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G15gat), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(G1gat), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g292(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT15), .B1(new_n470), .B2(new_n472), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n473), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n467), .A4(new_n464), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT17), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n504));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n507));
  AND4_X1   g306(.A1(new_n507), .A2(new_n482), .A3(new_n498), .A4(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n495), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT89), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n512), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n499), .B(KEYINPUT90), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n507), .B1(new_n502), .B2(KEYINPUT17), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n508), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n517), .B(new_n514), .C1(new_n519), .C2(new_n495), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT18), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n502), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n523), .B2(new_n495), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n514), .B(KEYINPUT13), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n521), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT11), .B(G169gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G197gat), .ZN(new_n531));
  XOR2_X1   g330(.A(G113gat), .B(G141gat), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT12), .Z(new_n534));
  NOR3_X1   g333(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n515), .A2(new_n522), .A3(KEYINPUT92), .A4(new_n526), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT93), .A3(new_n534), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT93), .B1(new_n540), .B2(new_n534), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n458), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  OR2_X1    g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  XOR2_X1   g346(.A(G57gat), .B(G64gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT94), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n546), .B1(new_n547), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n548), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT95), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n511), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n301), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G211gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n564), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n568), .B(new_n571), .Z(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT7), .ZN(new_n574));
  INV_X1    g373(.A(G99gat), .ZN(new_n575));
  INV_X1    g374(.A(G106gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT8), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n574), .B(new_n577), .C1(G85gat), .C2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT97), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n510), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT41), .ZN(new_n586));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  OAI221_X1 g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .C1(new_n502), .C2(new_n584), .ZN(new_n588));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT98), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n586), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n590), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n584), .A2(new_n555), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n559), .A3(new_n583), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT99), .A3(new_n600), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n584), .A2(KEYINPUT99), .A3(new_n555), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT10), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n601), .A2(G230gat), .A3(G233gat), .A4(new_n602), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(new_n311), .ZN(new_n609));
  INV_X1    g408(.A(G204gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT100), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n603), .B2(new_n605), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n615), .A2(new_n607), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n613), .B1(new_n616), .B2(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(new_n613), .C1(new_n616), .C2(new_n612), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n597), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n545), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(new_n364), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT102), .B(G1gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1324gat));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G8gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT104), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n545), .A2(new_n622), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n448), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n623), .A2(KEYINPUT103), .A3(new_n447), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n628), .A2(KEYINPUT104), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n628), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n631), .A2(KEYINPUT42), .A3(new_n448), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT105), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n632), .A2(new_n633), .A3(new_n285), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(G1325gat));
  NOR2_X1   g440(.A1(new_n450), .A2(new_n451), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n488), .B1(new_n623), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n444), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G15gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT106), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n623), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n623), .A2(new_n416), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n458), .A2(new_n595), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n527), .A2(new_n537), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n539), .A2(new_n528), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n534), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n535), .B1(new_n657), .B2(new_n541), .ZN(new_n658));
  NOR4_X1   g457(.A1(new_n652), .A2(new_n658), .A3(new_n572), .A4(new_n621), .ZN(new_n659));
  INV_X1    g458(.A(new_n364), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n460), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n544), .A2(KEYINPUT108), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n621), .A2(new_n572), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n595), .B(KEYINPUT109), .Z(new_n669));
  AND3_X1   g468(.A1(new_n458), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n458), .B2(new_n595), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n666), .B(new_n667), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n364), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n662), .A2(new_n673), .ZN(G1328gat));
  AND3_X1   g473(.A1(new_n659), .A2(new_n461), .A3(new_n448), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n672), .B2(new_n447), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(G1329gat));
  OAI21_X1  g479(.A(G43gat), .B1(new_n672), .B2(new_n444), .ZN(new_n681));
  INV_X1    g480(.A(new_n642), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n659), .A2(new_n471), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n672), .B2(new_n416), .ZN(new_n687));
  INV_X1    g486(.A(new_n416), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n659), .A2(new_n469), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n666), .A2(new_n597), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n458), .A2(new_n621), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n660), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n448), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT49), .ZN(new_n698));
  INV_X1    g497(.A(G64gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR3_X1    g499(.A1(new_n697), .A2(KEYINPUT110), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT110), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1333gat));
  AND2_X1   g504(.A1(new_n694), .A2(new_n682), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G71gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n694), .A2(G71gat), .A3(new_n644), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT50), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n707), .B(new_n714), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n694), .A2(new_n688), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT112), .B(G78gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1335gat));
  INV_X1    g518(.A(new_n621), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G85gat), .A3(new_n364), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT114), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n666), .A2(new_n572), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT51), .B1(new_n652), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n458), .A2(new_n726), .A3(new_n595), .A4(new_n723), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(KEYINPUT113), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT113), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n621), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n670), .B2(new_n671), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n364), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n733), .B2(new_n447), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n720), .A2(G92gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n725), .A2(new_n448), .A3(new_n727), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(KEYINPUT115), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n733), .B2(new_n444), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n575), .B(new_n621), .C1(new_n728), .C2(new_n729), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n642), .ZN(G1338gat));
  NAND2_X1  g542(.A1(new_n652), .A2(KEYINPUT44), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n458), .A2(new_n668), .A3(new_n669), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n731), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n576), .B1(new_n746), .B2(new_n688), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT53), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n688), .B(new_n732), .C1(new_n670), .C2(new_n671), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n621), .A2(new_n576), .A3(new_n688), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT116), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n725), .A2(new_n727), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n751), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n755), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT118), .B1(new_n747), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n751), .B2(KEYINPUT117), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(new_n764), .ZN(G1339gat));
  NAND2_X1  g564(.A1(new_n416), .A2(new_n455), .ZN(new_n766));
  INV_X1    g565(.A(new_n572), .ZN(new_n767));
  INV_X1    g566(.A(new_n613), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n603), .A2(new_n614), .A3(new_n605), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT54), .A3(new_n606), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n614), .C1(new_n603), .C2(new_n605), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n611), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n769), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n774), .A3(new_n769), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n768), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n657), .A2(new_n541), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n664), .B1(new_n779), .B2(new_n536), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT108), .B(new_n535), .C1(new_n657), .C2(new_n541), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n512), .A2(new_n514), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT119), .Z(new_n784));
  NOR2_X1   g583(.A1(new_n524), .A2(new_n525), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n533), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(new_n536), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n618), .A2(new_n787), .A3(new_n620), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n669), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n669), .A2(new_n778), .A3(new_n787), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n767), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n666), .A2(new_n597), .A3(new_n621), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n766), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n448), .A2(new_n364), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n218), .A3(new_n666), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n452), .B1(new_n792), .B2(new_n794), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n796), .ZN(new_n801));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n658), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(G1340gat));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n216), .A3(new_n621), .ZN(new_n804));
  OAI21_X1  g603(.A(G120gat), .B1(new_n801), .B2(new_n720), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n797), .B2(new_n767), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n795), .A2(KEYINPUT121), .A3(new_n572), .A4(new_n796), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n221), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n800), .A2(G127gat), .A3(new_n572), .A4(new_n796), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(KEYINPUT120), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(KEYINPUT120), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(G1342gat));
  OR4_X1    g613(.A1(KEYINPUT56), .A2(new_n797), .A3(G134gat), .A4(new_n596), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n228), .A3(new_n595), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n801), .B2(new_n596), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(G1343gat));
  INV_X1    g618(.A(new_n796), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n644), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n771), .A2(new_n774), .A3(new_n769), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n613), .B1(new_n823), .B2(new_n775), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n788), .B1(new_n824), .B2(new_n658), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n596), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n572), .B1(new_n826), .B2(new_n790), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n688), .B1(new_n827), .B2(new_n793), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n822), .B1(new_n828), .B2(KEYINPUT57), .ZN(new_n829));
  INV_X1    g628(.A(new_n669), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n663), .B2(new_n665), .ZN(new_n831));
  INV_X1    g630(.A(new_n788), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n572), .B1(new_n833), .B2(new_n790), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n688), .B1(new_n834), .B2(new_n793), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(KEYINPUT57), .ZN(new_n836));
  OAI21_X1  g635(.A(G141gat), .B1(new_n836), .B2(new_n658), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n822), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n658), .A2(G141gat), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n829), .B(new_n666), .C1(new_n835), .C2(KEYINPUT57), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n842), .A2(G141gat), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(G1344gat));
  AOI21_X1  g644(.A(new_n416), .B1(new_n792), .B2(new_n794), .ZN(new_n846));
  INV_X1    g645(.A(G148gat), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n621), .A4(new_n821), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n778), .A2(KEYINPUT123), .A3(new_n595), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n824), .B2(new_n596), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n856), .A3(new_n787), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n572), .B1(new_n857), .B2(new_n826), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n597), .A2(new_n544), .A3(new_n621), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n853), .B(new_n688), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n852), .A2(new_n621), .A3(new_n821), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n851), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n829), .B(new_n621), .C1(new_n835), .C2(KEYINPUT57), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(new_n851), .A3(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n850), .B1(new_n862), .B2(new_n864), .ZN(G1345gat));
  AOI21_X1  g664(.A(G155gat), .B1(new_n838), .B2(new_n572), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n836), .A2(new_n204), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n572), .ZN(G1346gat));
  AOI21_X1  g667(.A(G162gat), .B1(new_n838), .B2(new_n595), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n836), .A2(new_n205), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n669), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n660), .A2(new_n447), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n795), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n666), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n310), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n452), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n872), .C1(new_n834), .C2(new_n793), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(G169gat), .A3(new_n544), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1348gat));
  NOR3_X1   g683(.A1(new_n877), .A2(new_n311), .A3(new_n720), .ZN(new_n885));
  INV_X1    g684(.A(new_n873), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n621), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n311), .ZN(G1349gat));
  OAI21_X1  g687(.A(G183gat), .B1(new_n877), .B2(new_n767), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n572), .A2(new_n300), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n873), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT60), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n889), .B(new_n893), .C1(new_n873), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1350gat));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n595), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G190gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n886), .A2(new_n296), .A3(new_n669), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND2_X1  g701(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n896), .A2(G190gat), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(G1351gat));
  INV_X1    g704(.A(new_n872), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n644), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n860), .B(new_n907), .C1(new_n846), .C2(new_n853), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n658), .ZN(new_n909));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n835), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n666), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1352gat));
  NOR4_X1   g713(.A1(new_n835), .A2(G204gat), .A3(new_n720), .A4(new_n910), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n852), .A2(new_n621), .A3(new_n860), .ZN(new_n918));
  OAI21_X1  g717(.A(G204gat), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n916), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(G1353gat));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  OAI211_X1 g722(.A(G211gat), .B(new_n923), .C1(new_n908), .C2(new_n767), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n289), .A3(new_n572), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n852), .A2(new_n572), .A3(new_n860), .A4(new_n907), .ZN(new_n928));
  INV_X1    g727(.A(new_n925), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n928), .A2(G211gat), .A3(new_n929), .A4(new_n923), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n908), .B2(new_n596), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n290), .A3(new_n669), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


