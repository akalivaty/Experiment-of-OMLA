//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n470), .B2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n462), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(G2104), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(new_n479), .ZN(G160));
  NAND3_X1  g055(.A1(new_n472), .A2(G2105), .A3(new_n474), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(new_n475), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n484), .A2(new_n489), .ZN(G162));
  AND2_X1   g065(.A1(new_n472), .A2(new_n474), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G126), .A4(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT72), .B1(new_n481), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n472), .A2(new_n474), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n462), .A2(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(new_n463), .C1(new_n503), .C2(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n517), .A2(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n512), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n520), .A2(new_n519), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n516), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n511), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n517), .A2(new_n539), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  OAI211_X1 g118(.A(G43), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n523), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(G56), .B1(new_n520), .B2(new_n519), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n511), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  XNOR2_X1  g130(.A(new_n509), .B(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(G78), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n517), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n517), .B2(new_n561), .ZN(new_n563));
  OR2_X1    g138(.A1(KEYINPUT5), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(KEYINPUT5), .A2(G543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(new_n514), .B2(new_n515), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n560), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n517), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n566), .A2(G87), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(G288));
  INV_X1    g151(.A(G73), .ZN(new_n577));
  INV_X1    g152(.A(G543), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT76), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT76), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n532), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n578), .B1(new_n514), .B2(new_n515), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n523), .ZN(G305));
  AOI22_X1  g161(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n511), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n517), .A2(new_n589), .B1(new_n523), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n583), .A2(G54), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n516), .A2(new_n509), .A3(G92), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n556), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n481), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT78), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n488), .B2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n470), .A2(new_n468), .A3(G2105), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT13), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT83), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT84), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(G23), .ZN(new_n693));
  INV_X1    g268(.A(new_n574), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n689), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT33), .B(G1976), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n688), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n488), .A2(G131), .ZN(new_n704));
  OR2_X1    g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n706));
  INV_X1    g281(.A(G119), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n481), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  AOI21_X1  g287(.A(new_n689), .B1(G290), .B2(KEYINPUT86), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT86), .B2(G290), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n689), .A2(G24), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT85), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n712), .B(new_n718), .C1(new_n698), .C2(new_n699), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n701), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT89), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n702), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n702), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G2090), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT98), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n689), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n689), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G1966), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n606), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G4), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G160), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n734), .A2(new_n735), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n732), .B(new_n743), .C1(new_n742), .C2(new_n741), .ZN(new_n744));
  NOR2_X1   g319(.A1(G27), .A2(G29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G164), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G2078), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n702), .A2(G32), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G105), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n478), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G129), .B2(new_n482), .ZN(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n475), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n759), .B2(new_n702), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n689), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT99), .B(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n702), .B1(new_n768), .B2(G28), .ZN(new_n770));
  AND2_X1   g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NOR2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(G301), .A2(G16), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n689), .A2(G5), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n550), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n730), .A2(G1966), .ZN(new_n782));
  INV_X1    g357(.A(new_n776), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G1961), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n767), .A2(new_n778), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n744), .A2(new_n747), .A3(new_n762), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n734), .A2(new_n735), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n626), .A2(new_n702), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(KEYINPUT97), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(KEYINPUT97), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n702), .A2(G33), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  INV_X1    g369(.A(G139), .ZN(new_n795));
  OAI221_X1 g370(.A(new_n793), .B1(new_n794), .B2(new_n462), .C1(new_n475), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n702), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT93), .B(G2072), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n702), .A2(G26), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT28), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G116), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n482), .B2(G128), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n488), .A2(new_n807), .A3(G140), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n488), .B2(G140), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n811), .B2(new_n702), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT91), .B(G2067), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n790), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n726), .A2(G2090), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n728), .A2(new_n786), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n723), .A2(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  XOR2_X1   g394(.A(KEYINPUT103), .B(G860), .Z(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n606), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n516), .A2(new_n509), .A3(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(G67), .B1(new_n520), .B2(new_n519), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n511), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n825), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n564), .B2(new_n565), .ZN(new_n833));
  INV_X1    g408(.A(new_n828), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n830), .B(G651), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n546), .A2(new_n549), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n824), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n834), .B1(new_n509), .B2(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT100), .B1(new_n840), .B2(new_n511), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n566), .A2(G93), .B1(new_n583), .B2(G55), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n843), .A2(KEYINPUT102), .A3(new_n550), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT101), .B1(new_n843), .B2(new_n550), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n839), .A2(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n823), .B(new_n847), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n821), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(KEYINPUT39), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n843), .A2(new_n821), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n810), .A2(new_n507), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n810), .A2(new_n507), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n759), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n758), .A3(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n797), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n866));
  OR2_X1    g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n868), .B1(new_n475), .B2(new_n869), .C1(new_n870), .C2(new_n481), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n704), .B2(new_n708), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n709), .A2(new_n871), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n873), .A2(new_n631), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n631), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n874), .ZN(new_n878));
  INV_X1    g453(.A(new_n631), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n873), .A2(new_n631), .A3(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n797), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT106), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n858), .B(new_n860), .C1(new_n885), .C2(new_n863), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n865), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n865), .A2(new_n886), .ZN(new_n889));
  INV_X1    g464(.A(new_n883), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n484), .A2(new_n489), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n626), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n484), .A2(new_n621), .A3(new_n489), .A4(new_n625), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n740), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n740), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n895), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n880), .A2(new_n881), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n889), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n906), .A3(new_n887), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n906), .B1(new_n892), .B2(new_n893), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT40), .B1(new_n915), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G395));
  XOR2_X1   g496(.A(G303), .B(new_n574), .Z(new_n922));
  XNOR2_X1  g497(.A(G305), .B(new_n592), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n922), .B(new_n923), .Z(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n847), .B(new_n615), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n560), .A2(new_n600), .A3(new_n604), .A4(new_n567), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n560), .A2(new_n567), .B1(new_n600), .B2(new_n604), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(new_n605), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .A3(new_n927), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n926), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n925), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n925), .A3(new_n937), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n924), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  INV_X1    g517(.A(new_n924), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n942), .A2(new_n943), .A3(new_n938), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n837), .A2(G868), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(G295));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n945), .A2(new_n949), .A3(new_n947), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n945), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n550), .B1(new_n831), .B2(new_n836), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n829), .A2(new_n830), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n826), .A2(new_n825), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(new_n838), .A3(new_n824), .A4(new_n835), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT102), .B1(new_n843), .B2(new_n550), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n958), .A2(G301), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G301), .B1(new_n958), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G286), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n847), .A2(G171), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n958), .A2(G301), .A3(new_n964), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G168), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n967), .A2(new_n930), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n936), .B1(new_n967), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n953), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n970), .A3(new_n930), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n943), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n973), .A2(KEYINPUT112), .A3(new_n943), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n975), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n924), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT43), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n924), .B1(new_n971), .B2(new_n972), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n912), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n984), .B(new_n986), .C1(new_n978), .C2(new_n979), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT44), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n980), .B2(new_n982), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT43), .B(new_n986), .C1(new_n978), .C2(new_n979), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n758), .B(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G2067), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n810), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n709), .B(new_n711), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n592), .B(G1986), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n467), .A2(new_n1003), .A3(new_n479), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n496), .B2(new_n506), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1010), .B(G1384), .C1(new_n496), .C2(new_n506), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1009), .A2(new_n1011), .A3(G2078), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT53), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n507), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1004), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n777), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1012), .A2(KEYINPUT53), .ZN(new_n1022));
  OAI21_X1  g597(.A(G171), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(G301), .A3(new_n1020), .A4(new_n1013), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(G171), .B2(KEYINPUT127), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1015), .A2(new_n1005), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(G86), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n566), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n584), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT116), .B(new_n1034), .C1(new_n1035), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT116), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT49), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n694), .A2(G1976), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1033), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1006), .A2(new_n1004), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(G8), .A3(new_n1044), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1043), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G1971), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT113), .B(G2090), .Z(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1019), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(G8), .B(new_n1058), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1060), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT118), .B(new_n1004), .C1(new_n1006), .C2(new_n1017), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1066), .A2(new_n1018), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1004), .B1(new_n1006), .B2(new_n1017), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1070), .A3(new_n1061), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1032), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1051), .B(new_n1064), .C1(new_n1072), .C2(new_n1058), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1016), .A2(new_n742), .A3(new_n1004), .A4(new_n1018), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G168), .A2(new_n1032), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT51), .B1(new_n1079), .B2(KEYINPUT126), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1032), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1079), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1081), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1082), .A2(new_n1079), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1080), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1030), .A2(new_n1074), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1048), .A2(G2067), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1019), .B2(new_n735), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n605), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n606), .B(new_n1091), .C1(new_n1019), .C2(new_n735), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1009), .A2(new_n1011), .A3(G1996), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1031), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n550), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1100));
  AND2_X1   g675(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1099), .A2(new_n1100), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1095), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1070), .A2(new_n1018), .A3(new_n1066), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(G1956), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1106), .A2(new_n1108), .B1(new_n1059), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G299), .A2(KEYINPUT121), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1107), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1059), .A2(new_n1109), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1105), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT123), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1122), .A2(new_n1124), .A3(new_n1128), .A4(new_n1125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1120), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1114), .B1(new_n1131), .B2(new_n1093), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1090), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1082), .A2(KEYINPUT119), .A3(G168), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT119), .B1(new_n1082), .B2(G168), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1058), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1136), .A2(new_n1064), .A3(new_n1051), .A4(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1073), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1088), .A2(KEYINPUT62), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1073), .A2(new_n1023), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1147), .B(new_n1080), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1064), .ZN(new_n1150));
  INV_X1    g725(.A(G288), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1043), .A2(new_n1045), .A3(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1035), .B(KEYINPUT117), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1150), .A2(new_n1051), .B1(new_n1154), .B2(new_n1033), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1144), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1008), .B1(new_n1133), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1007), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1000), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1158), .A2(G1986), .A3(G290), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(KEYINPUT48), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(KEYINPUT48), .B2(new_n1160), .ZN(new_n1162));
  INV_X1    g737(.A(new_n997), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1007), .B1(new_n1163), .B2(new_n758), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1158), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1007), .B2(new_n994), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n709), .A2(new_n711), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n998), .A2(new_n1170), .B1(G2067), .B2(new_n810), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1007), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1162), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1157), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g749(.A1(new_n990), .A2(new_n991), .ZN(new_n1176));
  NOR4_X1   g750(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1177));
  AOI21_X1  g751(.A(KEYINPUT109), .B1(new_n908), .B2(new_n914), .ZN(new_n1178));
  NOR3_X1   g752(.A1(new_n917), .A2(new_n916), .A3(new_n913), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1176), .A2(new_n1180), .ZN(G308));
  OAI221_X1 g755(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .C1(new_n990), .C2(new_n991), .ZN(G225));
endmodule


