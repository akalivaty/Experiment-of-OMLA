//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  NAND2_X1  g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT93), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT92), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G57gat), .B(G64gat), .Z(new_n209));
  INV_X1    g008(.A(new_n203), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(KEYINPUT9), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n211), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT94), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(KEYINPUT94), .A3(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G127gat), .B(G155gat), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT20), .Z(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n222), .A2(new_n225), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n202), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n220), .B(new_n221), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n224), .ZN(new_n231));
  INV_X1    g030(.A(new_n202), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G1gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G1gat), .B2(new_n235), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G8gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n219), .B2(KEYINPUT21), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n242), .A3(new_n233), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(G162gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT8), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n256), .C1(G85gat), .C2(G92gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G99gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n263), .B2(new_n262), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT91), .B(G36gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G29gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT14), .ZN(new_n268));
  OR3_X1    g067(.A1(new_n268), .A2(G29gat), .A3(G36gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(G29gat), .B2(G36gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n265), .B1(new_n273), .B2(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n252), .B1(new_n260), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(KEYINPUT17), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n259), .B1(new_n275), .B2(KEYINPUT17), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n251), .B1(new_n281), .B2(KEYINPUT96), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(KEYINPUT97), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(KEYINPUT97), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n279), .B(new_n280), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n286), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n259), .B1(new_n217), .B2(new_n218), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n260), .A2(new_n215), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n259), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G120gat), .B(G148gat), .Z(new_n301));
  XNOR2_X1  g100(.A(G176gat), .B(G204gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n300), .B2(new_n303), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n305), .A3(new_n303), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n246), .A2(new_n290), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n239), .B1(new_n275), .B2(KEYINPUT17), .ZN(new_n312));
  INV_X1    g111(.A(new_n275), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n277), .A2(new_n312), .B1(new_n313), .B2(new_n239), .ZN(new_n314));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(KEYINPUT18), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n275), .B(new_n239), .Z(new_n317));
  XOR2_X1   g116(.A(new_n315), .B(KEYINPUT13), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT18), .B1(new_n314), .B2(new_n315), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G141gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(G197gat), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT11), .B(G169gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(KEYINPUT12), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n322), .B(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n311), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G1gat), .B(G29gat), .Z(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337));
  AND2_X1   g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(G113gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(G113gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n337), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n338), .A2(new_n339), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n345), .A2(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(G141gat), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n356), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G155gat), .B(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(G141gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(new_n362), .A3(new_n354), .A4(new_n356), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT82), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n352), .B1(new_n370), .B2(KEYINPUT1), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n349), .A2(new_n337), .A3(new_n372), .A4(new_n343), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n364), .A2(new_n371), .A3(new_n373), .A4(new_n368), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n369), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AND4_X1   g177(.A1(new_n354), .A2(new_n367), .A3(new_n362), .A4(new_n356), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT80), .B1(new_n365), .B2(new_n366), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n362), .B1(new_n380), .B2(new_n356), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n384), .A3(new_n368), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT81), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n379), .A2(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT5), .B1(new_n378), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n364), .A2(new_n368), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n383), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n369), .A2(new_n376), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n397), .B2(new_n388), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n394), .A3(new_n388), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n374), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n386), .B2(KEYINPUT4), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n377), .B1(new_n369), .B2(new_n376), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n388), .A2(KEYINPUT5), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n336), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n369), .A2(new_n376), .A3(new_n377), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n409), .A2(new_n389), .A3(new_n386), .A4(new_n391), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n397), .A2(new_n394), .A3(new_n388), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT5), .B(new_n410), .C1(new_n411), .C2(new_n398), .ZN(new_n412));
  INV_X1    g211(.A(new_n406), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n335), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n408), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416));
  OAI221_X1 g215(.A(new_n336), .B1(new_n416), .B2(KEYINPUT6), .C1(new_n401), .C2(new_n406), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  AND2_X1   g220(.A1(G211gat), .A2(G218gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(G211gat), .A2(G218gat), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT75), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G211gat), .ZN(new_n425));
  INV_X1    g224(.A(G218gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g227(.A1(G211gat), .A2(G218gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT22), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(KEYINPUT74), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G197gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G204gat), .ZN(new_n435));
  INV_X1    g234(.A(G204gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G197gat), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT74), .B1(new_n429), .B2(new_n432), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT76), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n424), .B(new_n430), .C1(new_n443), .C2(new_n439), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n440), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(KEYINPUT76), .A3(new_n424), .A4(new_n430), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(KEYINPUT29), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  INV_X1    g255(.A(G169gat), .ZN(new_n457));
  INV_X1    g256(.A(G176gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n459), .A2(KEYINPUT26), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463));
  NOR2_X1   g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n455), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT27), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G183gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G183gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT27), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n467), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n469), .A2(new_n475), .A3(KEYINPUT28), .A4(new_n472), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n474), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(G176gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n457), .A2(KEYINPUT64), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G169gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G169gat), .A2(G176gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT65), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n486), .B1(G169gat), .B2(G176gat), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n485), .A2(new_n491), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n460), .B2(new_n461), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n458), .A2(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT25), .B1(new_n500), .B2(G169gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(G183gat), .A2(G190gat), .ZN(new_n503));
  AND2_X1   g302(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(G190gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n455), .A2(new_n506), .A3(new_n481), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(new_n455), .B2(new_n481), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n480), .A2(new_n498), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n454), .B1(new_n479), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n459), .A2(KEYINPUT26), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n464), .A2(new_n456), .A3(new_n463), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n496), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n469), .A2(new_n475), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT67), .ZN(new_n516));
  AOI21_X1  g315(.A(G190gat), .B1(new_n469), .B2(new_n470), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT28), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n478), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n455), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n480), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n509), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT78), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n453), .B1(new_n511), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n477), .A2(new_n478), .ZN(new_n526));
  INV_X1    g325(.A(new_n466), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(new_n527), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n450), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n449), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n450), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n451), .A3(new_n524), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n448), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT79), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n531), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n421), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n531), .A2(new_n421), .A3(new_n536), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n536), .A4(new_n421), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n418), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n445), .A2(new_n447), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n384), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n395), .ZN(new_n552));
  NAND2_X1  g351(.A1(G228gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n385), .A2(new_n533), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n448), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n448), .A2(new_n554), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n532), .B1(new_n441), .B2(new_n444), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n395), .B1(new_n557), .B2(KEYINPUT3), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n552), .A2(new_n555), .B1(new_n559), .B2(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(G22gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT86), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G78gat), .B(G106gat), .Z(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G50gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n553), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n390), .B1(new_n550), .B2(new_n384), .ZN(new_n567));
  INV_X1    g366(.A(new_n553), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n566), .B(new_n561), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n567), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n568), .B1(new_n556), .B2(new_n558), .ZN(new_n572));
  OAI21_X1  g371(.A(G22gat), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n562), .A2(new_n565), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n575));
  AND4_X1   g374(.A1(new_n575), .A2(new_n573), .A3(new_n570), .A4(new_n565), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G227gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n383), .B1(new_n479), .B2(new_n510), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n520), .A2(new_n523), .A3(new_n581), .A4(new_n353), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n528), .B2(new_n353), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT32), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G15gat), .B(G43gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G99gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(KEYINPUT71), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT33), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n585), .B2(KEYINPUT32), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n587), .A2(new_n593), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n520), .A2(new_n523), .A3(new_n353), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT70), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n578), .A3(new_n582), .A4(new_n580), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT34), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n580), .A2(new_n582), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n578), .A4(new_n599), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n583), .A2(new_n584), .A3(new_n579), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT72), .B1(new_n607), .B2(new_n603), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n606), .B2(new_n608), .ZN(new_n612));
  INV_X1    g411(.A(new_n590), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n586), .A2(new_n596), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n585), .A2(KEYINPUT32), .A3(new_n593), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n607), .A2(KEYINPUT72), .A3(new_n603), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n604), .A2(new_n605), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT73), .A4(new_n601), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n577), .A2(new_n610), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT35), .B1(new_n548), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n548), .C2(new_n621), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n407), .A2(new_n408), .A3(new_n414), .ZN(new_n626));
  OAI211_X1 g425(.A(KEYINPUT6), .B(new_n336), .C1(new_n401), .C2(new_n406), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n577), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n618), .A3(new_n601), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n616), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n421), .ZN(new_n633));
  INV_X1    g432(.A(new_n540), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n539), .B1(new_n531), .B2(new_n536), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n544), .A4(new_n545), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n629), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n577), .A2(KEYINPUT87), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT87), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n574), .B2(new_n576), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n548), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n646), .B(new_n388), .C1(new_n403), .C2(new_n404), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n647), .A2(new_n335), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n369), .A2(new_n376), .A3(new_n389), .A4(new_n396), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT39), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT88), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n388), .B1(new_n403), .B2(new_n404), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT88), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n653), .A3(KEYINPUT39), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT40), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n335), .B1(new_n412), .B2(new_n413), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n648), .A2(KEYINPUT40), .A3(new_n655), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n659), .C1(new_n541), .C2(new_n546), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT37), .B1(new_n634), .B2(new_n635), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n531), .A2(new_n662), .A3(new_n536), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n663), .A2(KEYINPUT38), .A3(new_n633), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n448), .B1(new_n525), .B2(new_n530), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n534), .A2(new_n535), .A3(new_n449), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(KEYINPUT37), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n663), .A3(new_n633), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n661), .A2(new_n664), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n626), .A2(new_n542), .A3(new_n627), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n660), .B(new_n577), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT36), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n597), .A2(new_n609), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n616), .A2(new_n630), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n620), .A2(KEYINPUT36), .A3(new_n610), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n645), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n641), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n330), .A2(KEYINPUT99), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT99), .B1(new_n330), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n418), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(new_n547), .ZN(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n236), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  INV_X1    g491(.A(G8gat), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n684), .A2(new_n693), .A3(new_n688), .A4(new_n690), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n683), .A2(new_n547), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n692), .B(new_n694), .C1(KEYINPUT42), .C2(new_n695), .ZN(G1325gat));
  XOR2_X1   g495(.A(new_n678), .B(KEYINPUT101), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n683), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n632), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n683), .B2(new_n700), .ZN(G1326gat));
  AND2_X1   g500(.A1(new_n642), .A2(new_n644), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  AND3_X1   g504(.A1(new_n645), .A2(new_n672), .A3(new_n678), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n639), .B1(new_n622), .B2(new_n623), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n625), .ZN(new_n708));
  INV_X1    g507(.A(new_n290), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n244), .A2(new_n245), .ZN(new_n711));
  INV_X1    g510(.A(new_n329), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n712), .A3(new_n310), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n685), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n708), .B2(new_n709), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n680), .A2(KEYINPUT44), .A3(new_n290), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n713), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724), .B2(new_n418), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n718), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n719), .A2(new_n725), .A3(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n266), .B1(new_n728), .B2(KEYINPUT46), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n688), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n724), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n688), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n266), .B1(new_n734), .B2(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(new_n678), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n738), .A3(new_n713), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n632), .A2(G43gat), .ZN(new_n741));
  AND4_X1   g540(.A1(new_n680), .A2(new_n713), .A3(new_n290), .A4(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n722), .A3(new_n697), .A4(new_n713), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n742), .B1(new_n745), .B2(G43gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT47), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n744), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n744), .B(KEYINPUT107), .C1(new_n749), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1330gat));
  OAI21_X1  g556(.A(G50gat), .B1(new_n724), .B2(new_n577), .ZN(new_n758));
  INV_X1    g557(.A(G50gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n714), .A2(new_n759), .A3(new_n702), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(KEYINPUT48), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n760), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n733), .A2(new_n702), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G50gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g564(.A1(new_n711), .A2(new_n712), .A3(new_n709), .A4(new_n310), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n708), .A2(new_n766), .A3(KEYINPUT108), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT108), .B1(new_n708), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n418), .B(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g572(.A(new_n547), .B(KEYINPUT110), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  NOR2_X1   g579(.A1(new_n698), .A2(new_n205), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n767), .A2(new_n768), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT111), .Z(new_n783));
  OAI21_X1  g582(.A(new_n205), .B1(new_n769), .B2(new_n632), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT50), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n702), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g590(.A1(new_n246), .A2(new_n712), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n309), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n723), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G85gat), .B1(new_n794), .B2(new_n418), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n712), .A4(new_n246), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n680), .A2(new_n290), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n792), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT112), .B(new_n797), .C1(new_n798), .C2(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n310), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n418), .A2(G85gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n795), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  OAI21_X1  g604(.A(G92gat), .B1(new_n794), .B2(new_n547), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n796), .A2(new_n799), .A3(KEYINPUT113), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n775), .A2(new_n309), .A3(G92gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n797), .C1(new_n798), .C2(new_n792), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n723), .A2(new_n774), .A3(new_n793), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n814), .B2(G92gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n802), .A3(new_n808), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(G1337gat));
  XNOR2_X1  g619(.A(KEYINPUT115), .B(G99gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n794), .B2(new_n698), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n632), .A2(new_n821), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n803), .B2(new_n823), .ZN(G1338gat));
  OAI21_X1  g623(.A(G106gat), .B1(new_n794), .B2(new_n577), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n309), .A2(G106gat), .A3(new_n577), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n801), .A2(new_n802), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n723), .A2(new_n702), .A3(new_n793), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n807), .A2(new_n810), .A3(new_n827), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(KEYINPUT116), .A3(KEYINPUT53), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n833), .B2(KEYINPUT53), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(new_n771), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n296), .A2(new_n297), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n291), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n296), .A2(new_n292), .A3(new_n297), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n303), .B1(new_n298), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n307), .B2(new_n308), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n847), .B(new_n329), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n322), .A2(new_n328), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n314), .A2(new_n315), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n317), .A2(new_n318), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n326), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n309), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n290), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n849), .A2(new_n850), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n288), .B2(new_n289), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n847), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n246), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n311), .A2(new_n712), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n837), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n621), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(new_n775), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n346), .A3(new_n329), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n702), .A2(new_n632), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n418), .A3(new_n774), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n329), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT119), .B1(new_n872), .B2(G113gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(G1340gat));
  INV_X1    g674(.A(new_n870), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n774), .A2(new_n418), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n310), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G120gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n342), .A3(new_n310), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1341gat));
  INV_X1    g683(.A(new_n871), .ZN(new_n885));
  OAI21_X1  g684(.A(G127gat), .B1(new_n885), .B2(new_n246), .ZN(new_n886));
  INV_X1    g685(.A(G127gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n887), .A3(new_n711), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n709), .A2(new_n688), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n864), .A2(new_n890), .A3(new_n865), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT56), .Z(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n885), .B2(new_n709), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n577), .B1(new_n862), .B2(new_n863), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n678), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n859), .A2(new_n847), .A3(new_n860), .ZN(new_n900));
  INV_X1    g699(.A(new_n308), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n901), .A2(new_n306), .B1(new_n845), .B2(new_n844), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n329), .A2(new_n848), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n309), .A2(new_n856), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n709), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n711), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n246), .A2(new_n329), .A3(new_n290), .A4(new_n310), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n702), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n899), .B1(new_n908), .B2(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n909), .A3(new_n329), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G141gat), .ZN(new_n911));
  OR2_X1    g710(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n697), .A2(new_n577), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n712), .A2(G141gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n864), .A2(new_n775), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n911), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n911), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n864), .A2(new_n913), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n774), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n921), .B(G148gat), .C1(new_n923), .C2(new_n310), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n898), .A2(new_n909), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n925), .B2(new_n309), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n897), .B(new_n702), .C1(new_n906), .C2(new_n907), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n310), .B(new_n927), .C1(new_n896), .C2(new_n897), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n678), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n924), .B1(new_n930), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n925), .B2(new_n246), .ZN(new_n932));
  INV_X1    g731(.A(G155gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n933), .A3(new_n711), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n925), .B2(new_n709), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n891), .A2(new_n250), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n922), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n775), .A2(new_n621), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n868), .A2(new_n418), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n488), .A2(new_n490), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n685), .B1(new_n862), .B2(new_n863), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n939), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n941), .A2(new_n942), .A3(new_n329), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n771), .A2(new_n547), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n868), .A2(new_n869), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n329), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n950), .B2(G169gat), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT123), .B(new_n457), .C1(new_n949), .C2(new_n329), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(G1348gat));
  INV_X1    g752(.A(new_n949), .ZN(new_n954));
  OAI21_X1  g753(.A(G176gat), .B1(new_n954), .B2(new_n309), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n941), .A2(new_n458), .A3(new_n310), .A4(new_n945), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  AOI21_X1  g756(.A(new_n474), .B1(new_n949), .B2(new_n711), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n940), .A2(new_n515), .A3(new_n246), .ZN(new_n959));
  OR3_X1    g758(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT60), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT60), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1350gat));
  NOR2_X1   g761(.A1(new_n709), .A2(G190gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n945), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n868), .A2(new_n290), .A3(new_n869), .A4(new_n948), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n964), .B(KEYINPUT124), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1351gat));
  NOR3_X1   g772(.A1(new_n697), .A2(new_n577), .A3(new_n775), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n943), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n434), .B1(new_n975), .B2(new_n712), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n698), .A2(new_n948), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n927), .B(new_n978), .C1(new_n896), .C2(new_n897), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n329), .A2(G197gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(G1352gat));
  OAI21_X1  g781(.A(G204gat), .B1(new_n928), .B2(new_n977), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n309), .A2(G204gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n943), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n983), .A2(new_n987), .A3(new_n990), .A4(new_n986), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1353gat));
  OR2_X1    g791(.A1(new_n979), .A2(new_n246), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(G211gat), .B1(new_n979), .B2(new_n246), .ZN(new_n997));
  NAND2_X1  g796(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n943), .A2(new_n425), .A3(new_n711), .A4(new_n974), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n979), .B2(new_n709), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n943), .A2(new_n426), .A3(new_n290), .A4(new_n974), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(KEYINPUT127), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1003), .A2(new_n1007), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1006), .A2(new_n1008), .ZN(G1355gat));
endmodule


