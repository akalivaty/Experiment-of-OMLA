//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT64), .B(new_n207), .C1(new_n203), .C2(G137), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(G134), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT64), .B1(new_n210), .B2(new_n207), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n205), .B(new_n206), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n204), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(new_n203), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n215), .B1(new_n218), .B2(new_n208), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n214), .B1(new_n219), .B2(new_n206), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n213), .A2(new_n220), .B1(new_n206), .B2(new_n219), .ZN(new_n221));
  XNOR2_X1  g035(.A(G143), .B(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT0), .A3(G128), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n219), .A2(new_n214), .A3(new_n206), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n210), .A2(new_n204), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G146), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT1), .A3(G146), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n239), .B(new_n240), .C1(G128), .C2(new_n222), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n236), .A2(new_n238), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n233), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .A3(new_n240), .A4(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n230), .A2(new_n232), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n227), .A2(new_n248), .A3(KEYINPUT30), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n219), .A2(new_n206), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n228), .B2(new_n229), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(new_n225), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n221), .A2(KEYINPUT66), .A3(new_n226), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n232), .B(new_n241), .C1(new_n213), .C2(new_n220), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n230), .A2(KEYINPUT67), .A3(new_n232), .A4(new_n241), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n253), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n200), .B(new_n249), .C1(new_n259), .C2(KEYINPUT30), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n248), .B1(new_n252), .B2(new_n225), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n200), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT70), .A2(G237), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(G237), .ZN(new_n267));
  AOI21_X1  g081(.A(G953), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n276));
  NAND4_X1  g090(.A1(new_n260), .A2(new_n264), .A3(new_n273), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n261), .B2(new_n200), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n227), .A2(new_n248), .A3(KEYINPUT28), .A4(new_n263), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(new_n281), .C1(new_n259), .C2(new_n263), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n283));
  INV_X1    g097(.A(new_n273), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n278), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n284), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n275), .A4(new_n277), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT75), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n288), .B2(new_n294), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT32), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT78), .B(G902), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n263), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT76), .B1(new_n262), .B2(new_n263), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n264), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n308), .A2(KEYINPUT28), .B1(new_n309), .B2(new_n280), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n264), .A2(KEYINPUT77), .A3(new_n279), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n305), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n282), .A2(new_n284), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n260), .A2(new_n264), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT29), .B(new_n315), .C1(new_n316), .C2(new_n284), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n301), .A2(new_n303), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT9), .B(G234), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G221), .B1(new_n321), .B2(G902), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G140), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G227), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n323), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G104), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT83), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G104), .ZN(new_n331));
  INV_X1    g145(.A(G107), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G107), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n328), .A2(KEYINPUT3), .A3(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n334), .A2(new_n336), .A3(new_n340), .A4(new_n337), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(new_n343), .A3(G101), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n226), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n333), .B1(G104), .B2(new_n332), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n347), .A3(new_n241), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(KEYINPUT84), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT84), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n347), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT85), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n341), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n349), .B1(new_n243), .B2(new_n246), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT86), .A4(new_n357), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n363), .A3(new_n252), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n353), .A2(new_n363), .A3(KEYINPUT87), .A4(new_n252), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n327), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n353), .A2(new_n363), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n221), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n241), .B1(new_n355), .B2(new_n357), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n341), .A2(new_n347), .A3(new_n241), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n221), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n366), .B2(new_n367), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n371), .B(G469), .C1(new_n326), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(G469), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT87), .B1(new_n380), .B2(new_n252), .ZN(new_n381));
  INV_X1    g195(.A(new_n367), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n370), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n327), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT12), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n374), .B(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n326), .B(new_n386), .C1(new_n381), .C2(new_n382), .ZN(new_n387));
  AOI211_X1 g201(.A(G469), .B(new_n304), .C1(new_n384), .C2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n322), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(KEYINPUT70), .A2(G237), .ZN(new_n390));
  OAI211_X1 g204(.A(G214), .B(new_n324), .C1(new_n390), .C2(new_n265), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT70), .B(G237), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n394), .A2(KEYINPUT91), .A3(G214), .A4(new_n324), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n395), .A3(new_n237), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT92), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT92), .A4(new_n237), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n268), .A2(KEYINPUT93), .A3(G143), .A4(G214), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n391), .B2(new_n237), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT17), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n398), .B2(new_n399), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n206), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  INV_X1    g228(.A(G140), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G125), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(G146), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(G146), .B1(new_n413), .B2(new_n416), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n406), .A2(KEYINPUT17), .A3(G131), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n411), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n328), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n409), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n406), .A2(KEYINPUT18), .A3(G131), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n400), .A2(new_n425), .A3(new_n405), .A4(new_n426), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n412), .B(new_n235), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n424), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n409), .A2(new_n436), .A3(new_n206), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n435), .A2(new_n437), .A3(new_n427), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n412), .B(KEYINPUT19), .Z(new_n439));
  OAI21_X1  g253(.A(new_n417), .B1(new_n439), .B2(G146), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n407), .B2(new_n410), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n434), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n433), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G475), .ZN(new_n444));
  INV_X1    g258(.A(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n422), .A2(new_n424), .A3(new_n432), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n424), .B1(new_n422), .B2(new_n432), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G475), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n233), .A2(G143), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n233), .A2(G143), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n453), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT95), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n453), .C1(new_n454), .C2(KEYINPUT13), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n454), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n464), .A2(new_n453), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n203), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G116), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(G116), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n332), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(KEYINPUT96), .A3(G134), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n463), .A2(new_n466), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n193), .A3(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT97), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n475), .A3(new_n193), .A4(G122), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n468), .A2(new_n475), .ZN(new_n481));
  OAI21_X1  g295(.A(G107), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n332), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n465), .B(new_n203), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G217), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n321), .A2(new_n490), .A3(G953), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n474), .A2(new_n488), .A3(new_n491), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n305), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n495), .B2(new_n305), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G475), .B1(new_n433), .B2(new_n442), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT20), .A3(new_n445), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n448), .A2(new_n452), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(G234), .A2(G237), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n507), .A2(G952), .A3(new_n324), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n304), .A2(G953), .A3(new_n507), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT21), .B(G898), .Z(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT68), .B(G119), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT5), .B(new_n194), .C1(new_n515), .C2(new_n193), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n191), .A2(new_n517), .A3(G116), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(G113), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(new_n199), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n355), .A2(new_n357), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n199), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n354), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n354), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(G110), .B(G122), .Z(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT8), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n342), .A2(new_n200), .A3(new_n344), .ZN(new_n531));
  INV_X1    g345(.A(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n225), .A2(G125), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(G125), .B2(new_n241), .ZN(new_n535));
  INV_X1    g349(.A(G224), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT7), .B1(new_n536), .B2(G953), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n535), .B(new_n537), .Z(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n445), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n531), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n528), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT6), .A3(new_n533), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n536), .A2(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n535), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n548), .A3(new_n528), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n445), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G210), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n542), .A2(new_n550), .A3(new_n553), .A4(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G214), .B1(G237), .B2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT88), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n389), .A2(new_n514), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n515), .A2(new_n233), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT79), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT23), .B1(new_n515), .B2(new_n233), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n187), .A2(G128), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n565), .A2(new_n566), .B1(KEYINPUT23), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n191), .B2(G128), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT24), .B(G110), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n412), .A2(new_n235), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n417), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n568), .A2(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n420), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n324), .A2(G221), .A3(G234), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT80), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT22), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n201), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n581), .B2(new_n579), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n590), .A3(new_n305), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n490), .B1(new_n305), .B2(G234), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT25), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n596), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n590), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n319), .A2(new_n562), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(G472), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n295), .B2(new_n305), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(new_n602), .A3(new_n302), .ZN(new_n608));
  INV_X1    g422(.A(new_n389), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n555), .A2(KEYINPUT99), .A3(new_n556), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n552), .A2(new_n612), .A3(new_n554), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n611), .A2(new_n560), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n448), .A2(new_n452), .A3(new_n504), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n474), .A2(new_n488), .A3(new_n491), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n491), .B1(new_n474), .B2(new_n488), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n493), .A2(KEYINPUT33), .A3(new_n494), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n305), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G478), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n495), .A2(new_n496), .A3(new_n305), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n626), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g442(.A1(new_n513), .A2(new_n614), .A3(new_n615), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n610), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  XNOR2_X1  g446(.A(new_n513), .B(KEYINPUT101), .ZN(new_n633));
  INV_X1    g447(.A(new_n502), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n448), .A2(new_n452), .A3(new_n634), .A4(new_n504), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n614), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n610), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n607), .A2(new_n302), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(new_n582), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n599), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n598), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n562), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  OAI21_X1  g464(.A(new_n509), .B1(new_n511), .B2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n611), .A2(new_n560), .A3(new_n613), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n389), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n319), .A2(new_n654), .A3(new_n645), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n651), .B(KEYINPUT39), .Z(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n609), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n448), .A2(new_n452), .A3(new_n504), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n502), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n316), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n284), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n445), .B1(new_n308), .B2(new_n273), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n301), .A2(new_n303), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n557), .B(KEYINPUT38), .ZN(new_n672));
  INV_X1    g486(.A(new_n645), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n560), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n665), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n237), .ZN(G45));
  NAND3_X1  g490(.A1(new_n615), .A2(new_n628), .A3(new_n651), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n389), .A2(new_n653), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n319), .A2(new_n645), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  AOI22_X1  g494(.A1(new_n383), .A2(new_n327), .B1(new_n368), .B2(new_n386), .ZN(new_n681));
  OAI21_X1  g495(.A(G469), .B1(new_n681), .B2(new_n304), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n366), .A2(new_n367), .B1(new_n221), .B2(new_n369), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n387), .B1(new_n683), .B2(new_n326), .ZN(new_n684));
  INV_X1    g498(.A(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n305), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n322), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n319), .A2(new_n629), .A3(new_n603), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n319), .A2(new_n603), .A3(new_n637), .A4(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  AOI21_X1  g507(.A(new_n685), .B1(new_n684), .B2(new_n305), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n388), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n614), .A2(new_n695), .A3(KEYINPUT105), .A4(new_n322), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n687), .B2(new_n653), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n514), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n319), .A3(new_n700), .A4(new_n645), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR4_X1   g516(.A1(new_n687), .A2(new_n653), .A3(new_n502), .A4(new_n663), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n273), .B1(new_n310), .B2(new_n311), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n298), .B1(new_n704), .B2(new_n278), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n607), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n603), .A3(new_n707), .A4(new_n633), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  AOI21_X1  g523(.A(new_n304), .B1(new_n288), .B2(new_n294), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n645), .B(new_n705), .C1(new_n710), .C2(new_n606), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n677), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n699), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT106), .B(G125), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G27));
  AOI21_X1  g529(.A(KEYINPUT32), .B1(new_n295), .B2(new_n298), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n300), .B(new_n297), .C1(new_n288), .C2(new_n294), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n602), .B1(new_n718), .B2(new_n318), .ZN(new_n719));
  INV_X1    g533(.A(new_n677), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n560), .A2(new_n322), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n555), .A2(new_n556), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT107), .B1(new_n379), .B2(new_n388), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n686), .A2(new_n724), .A3(new_n378), .A4(new_n377), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n719), .A2(new_n720), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n319), .A2(new_n603), .A3(new_n720), .A4(new_n726), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  INV_X1    g550(.A(new_n652), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n319), .A2(new_n603), .A3(new_n737), .A4(new_n726), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  OAI21_X1  g553(.A(new_n371), .B1(new_n326), .B2(new_n376), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n371), .B(KEYINPUT45), .C1(new_n326), .C2(new_n376), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(G469), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n378), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT110), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n686), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n686), .C1(new_n745), .C2(new_n746), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(KEYINPUT110), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n322), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n657), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n625), .A2(new_n627), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n615), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(new_n641), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n645), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n557), .A2(new_n559), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n761), .A2(new_n762), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n756), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n754), .A2(new_n771), .A3(new_n322), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n754), .B2(new_n322), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n319), .A2(new_n603), .A3(new_n677), .A4(new_n765), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT112), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  NOR2_X1   g593(.A1(new_n670), .A2(new_n602), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n672), .A2(new_n615), .A3(new_n757), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n695), .B(KEYINPUT49), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n721), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AND4_X1   g597(.A1(KEYINPUT20), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT20), .B1(new_n503), .B2(new_n445), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n634), .A4(new_n452), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n635), .A2(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n615), .A2(new_n628), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n561), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n608), .A3(new_n609), .A4(new_n633), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n794), .A2(new_n604), .A3(new_n646), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n701), .A2(new_n692), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n689), .A2(new_n708), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT114), .B1(new_n506), .B2(new_n651), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  INV_X1    g614(.A(new_n651), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n505), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n379), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n722), .B1(new_n804), .B2(new_n686), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n319), .A2(new_n645), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n712), .A2(new_n726), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n738), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n735), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n798), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n653), .A2(new_n663), .A3(new_n502), .A4(new_n801), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n645), .B1(new_n723), .B2(new_n725), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n670), .A2(new_n322), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n655), .A3(new_n713), .A4(new_n679), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT53), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n689), .A2(new_n701), .A3(new_n692), .A4(new_n708), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n735), .A3(new_n795), .A4(new_n808), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n673), .B1(new_n718), .B2(new_n318), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n820), .A2(new_n654), .B1(new_n699), .B2(new_n712), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n815), .A3(new_n679), .A4(new_n813), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n695), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n722), .A3(new_n509), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n780), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n615), .A3(new_n628), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n687), .A2(KEYINPUT116), .A3(new_n560), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n672), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n607), .A2(new_n602), .A3(new_n706), .A4(new_n509), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n687), .B2(new_n560), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n759), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n837), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n759), .A2(new_n829), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(new_n711), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n773), .B2(new_n774), .ZN(new_n849));
  INV_X1    g663(.A(new_n774), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n772), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n828), .A2(new_n322), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n834), .A2(new_n759), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n765), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n847), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n856), .B1(new_n775), .B2(new_n852), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(KEYINPUT51), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n858), .A2(new_n859), .B1(new_n847), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n809), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n795), .A2(new_n797), .A3(new_n796), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n825), .B1(new_n819), .B2(new_n824), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(G952), .B(new_n324), .C1(new_n830), .C2(new_n790), .ZN(new_n869));
  INV_X1    g683(.A(new_n719), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n845), .A2(KEYINPUT48), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT48), .B1(new_n845), .B2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n834), .A2(new_n759), .A3(new_n699), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n827), .A2(new_n862), .A3(new_n868), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n783), .B1(new_n878), .B2(new_n879), .ZN(G75));
  OR2_X1    g694(.A1(new_n324), .A2(G952), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT121), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n305), .B1(new_n865), .B2(new_n866), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(new_n554), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n545), .A2(new_n549), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n547), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n887), .B(new_n888), .Z(new_n889));
  OR2_X1    g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n889), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(G51));
  XOR2_X1   g706(.A(new_n378), .B(KEYINPUT57), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n827), .B2(new_n868), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n895), .B2(new_n681), .ZN(new_n896));
  INV_X1    g710(.A(new_n744), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n865), .A2(new_n867), .A3(new_n866), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n684), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n896), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(new_n882), .ZN(G54));
  NAND3_X1  g719(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(new_n443), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n443), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n883), .B1(new_n907), .B2(new_n908), .ZN(G60));
  NAND2_X1  g723(.A1(new_n827), .A2(new_n868), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n619), .A2(new_n620), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n496), .A2(new_n445), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n915), .A2(KEYINPUT124), .A3(new_n882), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT124), .B1(new_n915), .B2(new_n882), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n911), .B1(new_n910), .B2(new_n914), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT60), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n865), .B2(new_n866), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(new_n643), .ZN(new_n923));
  INV_X1    g737(.A(new_n601), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n882), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n927), .B(KEYINPUT61), .C1(new_n923), .C2(new_n925), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G66));
  INV_X1    g746(.A(new_n512), .ZN(new_n933));
  OAI21_X1  g747(.A(G953), .B1(new_n933), .B2(new_n536), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n864), .B2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n886), .B1(G898), .B2(new_n324), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  OAI21_X1  g752(.A(new_n249), .B1(new_n259), .B2(KEYINPUT30), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n439), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n738), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n821), .A2(new_n679), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n768), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n719), .A2(new_n614), .A3(new_n664), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n756), .A2(new_n945), .B1(new_n734), .B2(new_n730), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n324), .A3(new_n778), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(G900), .A2(G953), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n659), .A2(new_n765), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n719), .A3(new_n791), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT127), .Z(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n675), .A2(new_n953), .A3(new_n943), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n675), .B2(new_n943), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n768), .B1(new_n775), .B2(new_n777), .ZN(new_n957));
  AOI211_X1 g771(.A(G953), .B(new_n940), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n324), .B1(G227), .B2(G900), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n949), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n947), .A2(new_n948), .ZN(new_n961));
  NAND2_X1  g775(.A1(G227), .A2(G900), .ZN(new_n962));
  AND4_X1   g776(.A1(G953), .A2(new_n961), .A3(new_n962), .A4(new_n940), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n944), .A2(new_n778), .A3(new_n946), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n798), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n316), .A2(new_n273), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n667), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n956), .A2(new_n864), .A3(new_n957), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n966), .ZN(new_n973));
  INV_X1    g787(.A(new_n969), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n966), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n667), .B(new_n975), .C1(new_n865), .C2(new_n866), .ZN(new_n976));
  NOR4_X1   g790(.A1(new_n970), .A2(new_n883), .A3(new_n973), .A4(new_n976), .ZN(G57));
endmodule


