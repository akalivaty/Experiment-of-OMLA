//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  OR2_X1    g0001(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OR2_X1    g0008(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(G50), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n211), .A2(new_n214), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G50), .A2(G226), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n216), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n219), .B(new_n230), .C1(new_n215), .C2(new_n218), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT14), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G232), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G226), .B2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G97), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n254), .A2(new_n259), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n251), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G238), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n249), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT13), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n265), .B(new_n270), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n247), .B1(new_n272), .B2(G169), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  AOI211_X1 g0074(.A(KEYINPUT14), .B(new_n274), .C1(new_n269), .C2(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  INV_X1    g0080(.A(G68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G20), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT12), .Z(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n212), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n248), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT72), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n255), .B2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(KEYINPUT69), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(G77), .B1(G50), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n293), .B2(G68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n286), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n284), .B(new_n290), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n278), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n272), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n269), .B2(new_n271), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n306), .A2(new_n302), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G238), .A2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n310), .B(new_n311), .C1(new_n252), .C2(G1698), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n264), .C1(G107), .C2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(new_n251), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n227), .C2(new_n267), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(G179), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  NOR2_X1   g0117(.A1(new_n255), .A2(G20), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT8), .A2(G58), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT8), .A2(G58), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n317), .A2(new_n318), .B1(new_n321), .B2(new_n296), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n293), .B2(new_n226), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n323), .A2(new_n286), .B1(new_n226), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n287), .A2(G77), .A3(new_n288), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n315), .A2(new_n274), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n316), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n304), .A2(new_n309), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n324), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n325), .B2(new_n286), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(new_n288), .ZN(new_n336));
  INV_X1    g0136(.A(G50), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n324), .A2(G50), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n342), .A2(G20), .A3(G33), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n295), .B2(new_n321), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(KEYINPUT70), .B(new_n343), .C1(new_n295), .C2(new_n321), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n293), .B1(new_n202), .B2(new_n203), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n339), .B(new_n341), .C1(new_n349), .C2(new_n287), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n295), .A2(new_n321), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT70), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  INV_X1    g0154(.A(new_n348), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n344), .A2(new_n345), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n340), .B1(new_n357), .B2(new_n286), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT9), .A3(new_n339), .ZN(new_n359));
  AND2_X1   g0159(.A1(KEYINPUT68), .A2(G223), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT68), .A2(G223), .ZN(new_n361));
  OAI21_X1  g0161(.A(G1698), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G222), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n310), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n264), .C1(G77), .C2(new_n310), .ZN(new_n366));
  INV_X1    g0166(.A(new_n267), .ZN(new_n367));
  INV_X1    g0167(.A(G226), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(KEYINPUT67), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n371), .A3(new_n314), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G200), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n305), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n352), .A2(new_n359), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n340), .B(new_n338), .C1(new_n357), .C2(new_n286), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n378), .B2(KEYINPUT9), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n373), .A4(new_n352), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n372), .A2(new_n274), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n372), .A2(G179), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n350), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n315), .A2(new_n305), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n315), .A2(G200), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n326), .A4(new_n327), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n257), .A2(KEYINPUT73), .A3(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n256), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n293), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n310), .B2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n281), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n281), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n207), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n296), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n391), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n293), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n410), .A3(new_n286), .ZN(new_n411));
  INV_X1    g0211(.A(new_n321), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n325), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n336), .B2(new_n412), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n368), .A2(G1698), .ZN(new_n416));
  OR2_X1    g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n310), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n251), .B1(new_n420), .B2(new_n264), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n267), .A2(new_n252), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT74), .B(G190), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n411), .A2(new_n415), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n404), .B1(new_n407), .B2(G68), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n287), .B1(new_n431), .B2(KEYINPUT16), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n414), .B1(new_n432), .B2(new_n405), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n425), .A4(new_n427), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n411), .A2(new_n415), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n274), .B1(new_n421), .B2(new_n423), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n263), .B1(new_n418), .B2(new_n419), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n437), .A2(new_n276), .A3(new_n422), .A4(new_n251), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT18), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n436), .A2(new_n438), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n433), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n430), .B(new_n434), .C1(new_n440), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n332), .A2(new_n387), .A3(new_n390), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G264), .A2(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(G257), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n310), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n257), .A2(G33), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n452));
  OAI21_X1  g0252(.A(G303), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT80), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT80), .B1(new_n450), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n264), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(G274), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n263), .ZN(new_n465));
  INV_X1    g0265(.A(G270), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n264), .C1(new_n454), .C2(new_n455), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n457), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n325), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n248), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n287), .A2(new_n324), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n293), .C1(G33), .C2(new_n260), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n286), .C1(new_n293), .C2(G116), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  OAI221_X1 g0284(.A(new_n476), .B1(new_n478), .B2(new_n475), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n474), .A2(G169), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n457), .A2(new_n471), .A3(new_n473), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(G179), .A4(new_n485), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n457), .A2(G179), .A3(new_n471), .A4(new_n473), .ZN(new_n492));
  INV_X1    g0292(.A(new_n485), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT82), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n474), .A2(KEYINPUT21), .A3(G169), .A4(new_n485), .ZN(new_n495));
  AND4_X1   g0295(.A1(new_n488), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n293), .B1(new_n255), .B2(new_n260), .ZN(new_n497));
  INV_X1    g0297(.A(G87), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n260), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(KEYINPUT19), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n256), .A2(new_n258), .A3(new_n293), .A4(G68), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n293), .A2(G33), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n260), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n286), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n212), .A2(new_n324), .A3(new_n285), .A4(new_n477), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n317), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n317), .A2(new_n324), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT77), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n310), .A2(new_n515), .A3(G244), .A4(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n310), .A2(G238), .A3(new_n363), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n264), .ZN(new_n520));
  INV_X1    g0320(.A(new_n460), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G250), .A3(new_n263), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n250), .B2(new_n521), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n512), .B1(new_n525), .B2(new_n274), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n519), .B2(new_n264), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n527), .A2(KEYINPUT78), .A3(new_n276), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT78), .B1(new_n527), .B2(new_n276), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n510), .B1(new_n506), .B2(new_n286), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n508), .A2(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n525), .B2(G200), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n305), .B2(new_n525), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n256), .A2(new_n258), .A3(new_n293), .A4(G87), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n310), .A2(KEYINPUT22), .A3(new_n293), .A4(G87), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n293), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n499), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n543), .B1(new_n318), .B2(G116), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT24), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n539), .A2(new_n540), .A3(new_n547), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n286), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n280), .A2(G20), .A3(new_n499), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n478), .A2(new_n499), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n287), .B1(new_n546), .B2(new_n548), .ZN(new_n557));
  INV_X1    g0357(.A(new_n555), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT83), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(G250), .A2(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n448), .A2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n256), .A2(new_n560), .A3(new_n258), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n458), .A2(new_n460), .B1(new_n213), .B2(new_n262), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n264), .A2(new_n564), .B1(new_n565), .B2(G264), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT84), .B1(new_n566), .B2(new_n461), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n264), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(G264), .ZN(new_n569));
  AND4_X1   g0369(.A1(KEYINPUT84), .A2(new_n568), .A3(new_n461), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G169), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(G179), .A3(new_n461), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n556), .A2(new_n559), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n550), .A2(new_n555), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(new_n461), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n461), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n305), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n307), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n536), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(new_n363), .ZN(new_n583));
  NOR2_X1   g0383(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n310), .A2(G250), .A3(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n479), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n583), .B2(new_n584), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT76), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n588), .ZN(new_n591));
  AND4_X1   g0391(.A1(G244), .A2(new_n256), .A3(new_n258), .A4(new_n363), .ZN(new_n592));
  INV_X1    g0392(.A(new_n584), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT76), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n583), .A2(new_n584), .B1(G33), .B2(G283), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n586), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n597), .A3(new_n264), .ZN(new_n598));
  INV_X1    g0398(.A(new_n461), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(G257), .B2(new_n565), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G169), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(G179), .A3(new_n600), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n324), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n499), .B1(new_n396), .B2(new_n398), .ZN(new_n605));
  INV_X1    g0405(.A(new_n296), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n226), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT6), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n260), .A2(new_n499), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G97), .A2(G107), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n499), .A2(KEYINPUT6), .A3(G97), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n293), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OR3_X1    g0413(.A1(new_n605), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n604), .B1(new_n614), .B2(new_n286), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n508), .A2(G97), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n602), .A2(new_n603), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n598), .A2(G190), .A3(new_n600), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n307), .B1(new_n598), .B2(new_n600), .ZN(new_n619));
  INV_X1    g0419(.A(new_n604), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n605), .A2(new_n607), .A3(new_n613), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n616), .C1(new_n621), .C2(new_n287), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n489), .A2(new_n426), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n493), .C1(new_n307), .C2(new_n489), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n496), .A2(new_n582), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n446), .A2(new_n627), .ZN(G372));
  NOR2_X1   g0428(.A1(new_n440), .A2(new_n443), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n278), .A2(new_n303), .B1(new_n309), .B2(new_n330), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n430), .A2(new_n434), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n382), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n385), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n623), .A2(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n520), .A2(KEYINPUT85), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n519), .A2(new_n639), .A3(new_n264), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n523), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT87), .B1(new_n641), .B2(new_n307), .ZN(new_n642));
  INV_X1    g0442(.A(new_n640), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n639), .B1(new_n519), .B2(new_n264), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n524), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G200), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n533), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n532), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n650), .B1(G190), .B2(new_n527), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n637), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n581), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n488), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n571), .A2(new_n572), .B1(new_n550), .B2(new_n555), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n617), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n658), .B2(new_n536), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT86), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n641), .B2(G169), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n645), .A2(KEYINPUT86), .A3(new_n274), .ZN(new_n663));
  INV_X1    g0463(.A(new_n512), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n527), .A2(new_n276), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n636), .B1(new_n446), .B2(new_n668), .ZN(G369));
  NOR2_X1   g0469(.A1(new_n573), .A2(new_n581), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n556), .A2(new_n559), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n279), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n248), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT89), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT91), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT91), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n670), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n496), .A2(new_n679), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n679), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n656), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n689), .A2(new_n493), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n655), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n496), .A2(new_n626), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(KEYINPUT90), .B(G330), .Z(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n573), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n685), .B1(new_n698), .B2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n217), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G1), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n500), .A2(G116), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n211), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(new_n689), .C1(new_n659), .C2(new_n667), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n666), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n652), .A2(new_n617), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(KEYINPUT26), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT26), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n617), .A2(new_n715), .A3(new_n530), .A4(new_n535), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT93), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(KEYINPUT26), .ZN(new_n718));
  AND4_X1   g0518(.A1(KEYINPUT93), .A2(new_n718), .A3(new_n666), .A4(new_n716), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n624), .B1(new_n655), .B2(new_n573), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n666), .A2(new_n654), .A3(new_n652), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n496), .A2(new_n698), .ZN(new_n725));
  INV_X1    g0525(.A(new_n723), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT94), .A4(new_n624), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n689), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n711), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  INV_X1    g0530(.A(new_n601), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n575), .A3(new_n474), .A4(new_n645), .ZN(new_n733));
  INV_X1    g0533(.A(new_n492), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT92), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(KEYINPUT30), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n527), .A2(new_n566), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n731), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n731), .A3(new_n738), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n736), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n733), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n679), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT31), .B(new_n743), .C1(new_n627), .C2(new_n679), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n745), .A3(new_n679), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n696), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n708), .B1(new_n749), .B2(G1), .ZN(G364));
  XNOR2_X1  g0550(.A(new_n697), .B(KEYINPUT95), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n705), .B1(G45), .B2(new_n672), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n751), .B(new_n753), .C1(new_n696), .C2(new_n695), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n212), .B1(G20), .B2(new_n274), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n276), .A2(G200), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(G20), .A3(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n498), .ZN(new_n760));
  NAND2_X1  g0560(.A1(G20), .A2(G179), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G200), .A3(new_n426), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n307), .A3(new_n426), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n337), .A2(new_n763), .B1(new_n764), .B2(new_n400), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n305), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n307), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n760), .B(new_n765), .C1(G68), .C2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n762), .A2(new_n305), .A3(new_n307), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G77), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n293), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n758), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G107), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n782), .A2(KEYINPUT32), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n293), .B1(new_n781), .B2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  OAI21_X1  g0587(.A(KEYINPUT32), .B1(new_n782), .B2(new_n783), .ZN(new_n788));
  AND4_X1   g0588(.A1(new_n310), .A2(new_n784), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n768), .A2(new_n776), .A3(new_n780), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n259), .B1(new_n791), .B2(new_n785), .C1(new_n759), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n763), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G326), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n769), .B1(new_n764), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n767), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G329), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n779), .A2(G283), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n795), .A2(new_n800), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n756), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n755), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n242), .A2(G45), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n702), .A2(new_n310), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(G45), .C2(new_n211), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n310), .A2(G355), .A3(new_n217), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G116), .C2(new_n217), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n805), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n808), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n695), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n754), .B1(new_n753), .B2(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n679), .A2(new_n328), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n390), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n330), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n331), .A2(new_n689), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n668), .B2(new_n679), .ZN(new_n824));
  INV_X1    g0624(.A(new_n823), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n689), .B(new_n825), .C1(new_n659), .C2(new_n667), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(new_n747), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n753), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n775), .A2(G116), .B1(G303), .B2(new_n794), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  INV_X1    g0631(.A(new_n767), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n779), .A2(G87), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n259), .B1(new_n796), .B2(new_n782), .C1(new_n764), .C2(new_n791), .ZN(new_n836));
  INV_X1    g0636(.A(new_n759), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G107), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g0638(.A1(new_n787), .A2(new_n834), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n764), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G137), .A2(new_n794), .B1(new_n840), .B2(G143), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n342), .B2(new_n832), .C1(new_n774), .C2(new_n783), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n310), .B1(new_n400), .B2(new_n785), .C1(new_n759), .C2(new_n337), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G68), .B2(new_n779), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n844), .B(new_n848), .C1(G132), .C2(new_n801), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n755), .B1(new_n839), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n755), .A2(new_n806), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n823), .A2(new_n806), .B1(new_n226), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(new_n752), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n829), .A2(new_n853), .ZN(G384));
  OAI21_X1  g0654(.A(new_n432), .B1(KEYINPUT16), .B2(new_n431), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n677), .B1(new_n855), .B2(new_n415), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n444), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n855), .A2(new_n415), .B1(new_n442), .B2(new_n677), .ZN(new_n858));
  INV_X1    g0658(.A(new_n428), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n677), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n435), .B1(new_n439), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n428), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n864));
  OAI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n857), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n435), .A2(new_n861), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n629), .B2(new_n631), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT107), .ZN(new_n870));
  INV_X1    g0670(.A(new_n864), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT106), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(new_n863), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT107), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n444), .A2(new_n875), .A3(new_n868), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n304), .A2(new_n689), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT105), .Z(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n857), .A2(new_n865), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n878), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n857), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n880), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n629), .A2(new_n677), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n822), .B(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n826), .A2(new_n896), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n302), .B(new_n679), .C1(new_n898), .C2(new_n309), .ZN(new_n899));
  INV_X1    g0699(.A(new_n309), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n302), .A2(new_n679), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n900), .B(new_n901), .C1(new_n278), .C2(new_n303), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n903), .ZN(new_n906));
  AOI211_X1 g0706(.A(KEYINPUT103), .B(new_n906), .C1(new_n826), .C2(new_n896), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n887), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n891), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n724), .A2(new_n727), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n718), .A2(new_n666), .A3(new_n716), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT93), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n714), .A2(KEYINPUT93), .A3(new_n716), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n679), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n710), .B1(new_n918), .B2(new_n709), .ZN(new_n919));
  INV_X1    g0719(.A(new_n446), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n635), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n911), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n823), .B1(new_n899), .B2(new_n902), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n744), .A2(new_n746), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n924), .B2(new_n879), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT40), .B1(new_n885), .B2(new_n886), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n926), .A2(new_n744), .A3(new_n746), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n744), .A2(new_n746), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n446), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n928), .B(new_n930), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n696), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n922), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n248), .B2(new_n672), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n611), .A2(new_n612), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT35), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n214), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(G116), .C1(new_n936), .C2(new_n935), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(G77), .B1(new_n400), .B2(new_n281), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n211), .A2(new_n940), .B1(G50), .B2(new_n281), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n279), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n939), .A3(new_n942), .ZN(G367));
  INV_X1    g0743(.A(KEYINPUT111), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n617), .A2(new_n679), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT108), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n679), .A2(new_n622), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n624), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n700), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n688), .B2(new_n951), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n698), .B1(new_n947), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n689), .B1(new_n956), .B2(new_n617), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n950), .A2(new_n686), .A3(new_n687), .A4(new_n953), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n679), .A2(new_n649), .A3(new_n650), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n666), .A2(new_n652), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n666), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n965), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n967), .A3(new_n963), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n952), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n944), .B1(new_n969), .B2(KEYINPUT110), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  INV_X1    g0771(.A(new_n952), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n967), .B1(new_n959), .B2(new_n963), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT111), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n970), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n974), .B1(new_n970), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n248), .B1(new_n672), .B2(G45), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n688), .A2(new_n690), .A3(new_n950), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT44), .B1(new_n691), .B2(new_n950), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n700), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n688), .B1(new_n699), .B2(new_n687), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n751), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n749), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT112), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n987), .A2(new_n749), .A3(new_n993), .A4(new_n990), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n748), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n703), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n981), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n980), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n837), .A2(G116), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT46), .Z(new_n1001));
  OAI22_X1  g0801(.A1(new_n832), .A2(new_n791), .B1(new_n796), .B2(new_n763), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n764), .A2(new_n792), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n259), .B1(new_n499), .B2(new_n785), .C1(new_n778), .C2(new_n260), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n831), .B2(new_n774), .C1(new_n1006), .C2(new_n782), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n782), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n310), .B1(new_n778), .B2(new_n226), .ZN(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n832), .A2(new_n783), .B1(new_n1011), .B2(new_n763), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G58), .C2(new_n837), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n786), .A2(G68), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n764), .B2(new_n342), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT113), .Z(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(new_n337), .C2(new_n774), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n753), .B1(new_n1019), .B2(new_n755), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n317), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n811), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n809), .B1(new_n217), .B2(new_n1021), .C1(new_n238), .C2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1020), .B(new_n1023), .C1(new_n962), .C2(new_n816), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n999), .A2(new_n1024), .ZN(G387));
  OAI22_X1  g0825(.A1(new_n774), .A2(new_n792), .B1(new_n1006), .B2(new_n764), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT114), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1026), .A2(new_n1027), .B1(new_n796), .B2(new_n832), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n797), .B2(new_n763), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n831), .B2(new_n785), .C1(new_n791), .C2(new_n759), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n801), .A2(G326), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n778), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n310), .B1(new_n1037), .B2(G116), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1021), .A2(new_n785), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n310), .B1(new_n782), .B2(new_n342), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n779), .C2(G97), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n767), .A2(new_n321), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G68), .A2(new_n770), .B1(new_n794), .B2(G159), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n837), .A2(G77), .B1(G50), .B2(new_n840), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n756), .B1(new_n1039), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n321), .A2(new_n337), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n706), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1049), .B(new_n459), .C1(KEYINPUT50), .C2(new_n1048), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G68), .B2(G77), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n811), .B1(new_n235), .B2(new_n459), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n706), .A2(new_n217), .A3(new_n310), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n217), .A2(G107), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n809), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n699), .B2(new_n816), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1047), .A2(new_n753), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n981), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n990), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n749), .A2(new_n990), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n749), .A2(new_n990), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n703), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(G393));
  XNOR2_X1  g0864(.A(new_n987), .B(new_n988), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n981), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n809), .B1(new_n260), .B2(new_n217), .C1(new_n245), .C2(new_n1022), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n782), .A2(new_n797), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n259), .B1(new_n475), .B2(new_n785), .C1(new_n759), .C2(new_n831), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G294), .B2(new_n770), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n796), .A2(new_n764), .B1(new_n763), .B2(new_n1006), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n767), .A2(G303), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n780), .A4(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n342), .A2(new_n763), .B1(new_n764), .B2(new_n783), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n835), .C1(new_n281), .C2(new_n759), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n786), .A2(G77), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n310), .B1(new_n782), .B2(new_n1011), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n767), .B2(G50), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n774), .C2(new_n412), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1068), .A2(new_n1074), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n753), .B1(new_n1082), .B2(new_n755), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1067), .B(new_n1083), .C1(new_n950), .C2(new_n816), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1066), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1065), .A2(new_n1062), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n992), .A2(new_n994), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n703), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(new_n879), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n894), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n918), .B2(new_n825), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n882), .B(new_n1092), .C1(new_n1094), .C2(new_n906), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n897), .A2(new_n903), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n882), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n880), .A2(new_n888), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n744), .A2(new_n923), .A3(new_n696), .A4(new_n746), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n744), .A2(G330), .A3(new_n746), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n923), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1059), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1098), .A2(new_n806), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n851), .A2(new_n412), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n259), .B1(new_n791), .B2(new_n782), .C1(new_n763), .C2(new_n831), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n779), .B2(G68), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n260), .B2(new_n774), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1078), .B1(new_n475), .B2(new_n764), .C1(new_n832), .C2(new_n499), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1112), .A2(new_n760), .A3(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT120), .Z(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n782), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n775), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n759), .A2(new_n342), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G128), .A2(new_n794), .B1(new_n840), .B2(G132), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n310), .B1(new_n783), .B2(new_n785), .C1(new_n778), .C2(new_n337), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G137), .B2(new_n767), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n753), .B1(new_n1127), .B2(new_n755), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1108), .A2(new_n1109), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1107), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n930), .A2(G330), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n636), .B(new_n1131), .C1(new_n730), .C2(new_n446), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT115), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n906), .B1(new_n747), .B2(new_n823), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1104), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n897), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT116), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n744), .A2(new_n1138), .A3(G330), .A4(new_n746), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n825), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n906), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n689), .B(new_n825), .C1(new_n720), .C2(new_n728), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1142), .A2(new_n894), .A3(new_n1100), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT117), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1136), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1105), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1133), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1096), .A2(new_n882), .B1(new_n880), .B2(new_n888), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1142), .A2(new_n894), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n879), .B1(new_n1151), .B2(new_n903), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1152), .B2(new_n882), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1153), .B2(new_n1104), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1136), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT117), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT117), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT115), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1132), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n921), .A2(KEYINPUT115), .A3(new_n1131), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1154), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1149), .A2(new_n1165), .A3(new_n703), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1149), .A2(new_n1165), .A3(KEYINPUT118), .A4(new_n703), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1130), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  NAND2_X1  g0971(.A1(new_n928), .A2(G330), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT124), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n386), .A2(KEYINPUT55), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT55), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n382), .A2(new_n1175), .A3(new_n385), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n378), .A2(new_n677), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1175), .B1(new_n382), .B2(new_n385), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n385), .ZN(new_n1181));
  AOI211_X1 g0981(.A(KEYINPUT55), .B(new_n1181), .C1(new_n377), .C2(new_n381), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1177), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1173), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1172), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n928), .A2(new_n1187), .A3(G330), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1189), .A2(new_n891), .A3(new_n910), .A4(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n928), .A2(G330), .A3(new_n1187), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1187), .B1(new_n928), .B2(G330), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n904), .A2(new_n907), .A3(new_n887), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n889), .A2(new_n890), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1192), .A2(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1059), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n806), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n832), .A2(new_n260), .B1(new_n1021), .B2(new_n769), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n259), .B1(new_n759), .B2(new_n226), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G41), .B1(new_n801), .B2(G283), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n778), .B2(new_n400), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1014), .B1(new_n763), .B2(new_n475), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n499), .C2(new_n764), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1116), .A2(new_n763), .B1(new_n769), .B2(new_n1008), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n837), .A2(new_n1118), .ZN(new_n1212));
  INV_X1    g1012(.A(G132), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1212), .B1(new_n342), .B2(new_n785), .C1(new_n1213), .C2(new_n832), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(G128), .C2(new_n840), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT59), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G41), .B1(new_n1037), .B2(G159), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G33), .B1(new_n801), .B2(G124), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n257), .A2(new_n255), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n337), .B1(new_n1221), .B2(G41), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1210), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1223), .A2(new_n755), .B1(new_n337), .B2(new_n851), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1199), .A2(new_n752), .A3(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1198), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1164), .B1(new_n1106), .B2(new_n1146), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT125), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1191), .A2(new_n1196), .A3(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n911), .B(KEYINPUT125), .C1(new_n1193), .C2(new_n1192), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(KEYINPUT57), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n703), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1133), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1197), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1232), .B2(new_n1234), .ZN(G375));
  NOR2_X1   g1035(.A1(new_n759), .A2(new_n783), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n259), .B(new_n1236), .C1(G128), .C2(new_n801), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n767), .A2(new_n1118), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1037), .A2(G58), .B1(G50), .B2(new_n786), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1213), .A2(new_n763), .B1(new_n769), .B2(new_n342), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G137), .B2(new_n840), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n259), .B1(new_n792), .B2(new_n782), .C1(new_n763), .C2(new_n791), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1040), .B(new_n1243), .C1(G97), .C2(new_n837), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n775), .A2(G107), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n779), .A2(G77), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n767), .A2(G116), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n764), .A2(new_n831), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1242), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1250), .A2(new_n755), .B1(new_n281), .B2(new_n851), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n752), .B(new_n1251), .C1(new_n903), .C2(new_n807), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1160), .B2(new_n981), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT126), .B(new_n1252), .C1(new_n1160), .C2(new_n981), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1133), .A2(new_n1146), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n996), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  INV_X1    g1061(.A(new_n1130), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1262), .A2(new_n1166), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G375), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(G384), .A3(G381), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n999), .A2(new_n1090), .A3(new_n1024), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1268), .A2(G396), .A3(G393), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(G407));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G343), .C2(new_n1266), .ZN(G409));
  AND3_X1   g1071(.A1(new_n1233), .A2(new_n996), .A3(new_n1197), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1229), .A2(new_n1059), .A3(new_n1230), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1225), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1262), .B(new_n1166), .C1(new_n1272), .C2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1170), .B2(G375), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1259), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1160), .A2(KEYINPUT60), .A3(new_n1164), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n703), .A3(new_n1258), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1257), .A2(new_n1280), .A3(G384), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1257), .B2(new_n1280), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n678), .A2(G213), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1276), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1276), .A2(new_n1285), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1283), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1281), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1287), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT63), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(G393), .B(G396), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1268), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1090), .B1(new_n999), .B2(new_n1024), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(G390), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1268), .A3(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1286), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1295), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1276), .A2(new_n1285), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT62), .B1(new_n1309), .B2(new_n1286), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1306), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1303), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1307), .A2(new_n1313), .ZN(G405));
  AND2_X1   g1114(.A1(G375), .A2(new_n1263), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1170), .A2(G375), .ZN(new_n1316));
  OR3_X1    g1116(.A1(new_n1284), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1284), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1317), .A2(new_n1318), .B1(new_n1303), .B2(KEYINPUT127), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1303), .B(KEYINPUT127), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(G402));
endmodule


