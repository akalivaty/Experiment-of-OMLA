//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT80), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n189), .B(new_n190), .Z(new_n191));
  XNOR2_X1  g005(.A(G104), .B(G107), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT81), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G107), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n193), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(G104), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(G101), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n194), .A2(new_n201), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(KEYINPUT64), .A3(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT64), .B1(new_n209), .B2(G143), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n206), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n222));
  AND4_X1   g036(.A1(KEYINPUT0), .A2(new_n210), .A3(new_n212), .A4(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n210), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(KEYINPUT64), .A3(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n220), .A2(new_n230), .A3(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT10), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n194), .A2(new_n201), .A3(new_n205), .ZN(new_n234));
  INV_X1    g048(.A(new_n213), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n236), .A2(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n219), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT67), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n246), .B2(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(G134), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n249), .ZN(new_n254));
  AOI211_X1 g068(.A(new_n243), .B(new_n248), .C1(new_n251), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n254), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n245), .A2(new_n247), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n242), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n241), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n253), .B1(new_n252), .B2(new_n249), .ZN(new_n260));
  AOI211_X1 g074(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n244), .C2(G134), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n243), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n248), .B1(new_n251), .B2(new_n254), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n242), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n240), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n259), .A2(new_n266), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n219), .A2(new_n232), .A3(new_n239), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n191), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n191), .B1(new_n240), .B2(new_n267), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n213), .B1(new_n217), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(new_n201), .A3(new_n205), .A4(new_n194), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n206), .B2(new_n218), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n259), .A3(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n263), .B2(new_n265), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n278), .A2(new_n279), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n273), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n279), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n280), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n284), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n272), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G469), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n191), .B1(new_n281), .B2(new_n271), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n269), .A2(new_n270), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(G469), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G469), .A2(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G221), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(new_n289), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT79), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT83), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n296), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n259), .A2(new_n229), .A3(new_n266), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n252), .B2(new_n247), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n264), .B2(new_n309), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n218), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n319), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n314), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n229), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n274), .A2(KEYINPUT0), .A3(G128), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n216), .B2(new_n227), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n263), .A2(new_n265), .B1(new_n328), .B2(KEYINPUT65), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n257), .B(new_n309), .C1(new_n260), .C2(new_n261), .ZN(new_n330));
  INV_X1    g144(.A(new_n310), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n217), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n235), .B1(new_n226), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT68), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n311), .A2(new_n336), .A3(new_n218), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n326), .A2(new_n329), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n313), .B(new_n324), .C1(new_n338), .C2(KEYINPUT30), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n324), .B(KEYINPUT70), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n308), .A2(new_n312), .A3(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G210), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n342), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G101), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n339), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT31), .ZN(new_n349));
  INV_X1    g163(.A(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n335), .A2(new_n337), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n328), .A2(KEYINPUT65), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n326), .C1(new_n258), .C2(new_n255), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n324), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n351), .B1(new_n356), .B2(new_n341), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n341), .A2(new_n351), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT31), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n339), .A2(new_n360), .A3(new_n341), .A4(new_n347), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n349), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(G472), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n357), .A2(new_n358), .A3(new_n350), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n347), .B1(new_n339), .B2(new_n341), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n368), .A2(KEYINPUT29), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n308), .A2(new_n312), .ZN(new_n371));
  INV_X1    g185(.A(new_n340), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n341), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n358), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n350), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n289), .ZN(new_n379));
  OAI21_X1  g193(.A(G472), .B1(new_n370), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n362), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  OR3_X1    g199(.A1(new_n385), .A2(KEYINPUT16), .A3(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(G146), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n209), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT75), .ZN(new_n392));
  INV_X1    g206(.A(G110), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT24), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G110), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G119), .B(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n207), .A2(G119), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n316), .A2(G128), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT24), .B(G110), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT75), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n316), .A2(G128), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT74), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT23), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n406), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(KEYINPUT23), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n411), .A2(new_n393), .A3(new_n401), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n391), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n414), .A2(new_n391), .A3(new_n404), .A4(new_n399), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n390), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n384), .A2(new_n386), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n209), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n387), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n401), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(KEYINPUT74), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n400), .B1(new_n412), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI221_X1 g239(.A(new_n421), .B1(new_n402), .B2(new_n403), .C1(new_n425), .C2(new_n393), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G137), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n422), .A2(new_n424), .A3(G110), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n399), .A2(new_n404), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT76), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n389), .B1(new_n434), .B2(new_n416), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n420), .A2(new_n387), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n425), .A2(new_n393), .B1(new_n402), .B2(new_n403), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n429), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n439), .A3(new_n289), .ZN(new_n440));
  NOR2_X1   g254(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(G217), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(G217), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(G234), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT73), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n431), .A2(new_n439), .A3(new_n289), .A4(new_n441), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n447), .A2(G902), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n431), .A2(new_n439), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT78), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G122), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G113), .B1(new_n317), .B2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n457), .A2(new_n459), .B1(new_n315), .B2(new_n320), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n206), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n222), .A2(new_n324), .A3(new_n231), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n462), .A3(new_n455), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(KEYINPUT6), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n328), .A2(G125), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n334), .A2(new_n385), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G224), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G953), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT85), .B(KEYINPUT6), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n463), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n463), .B2(new_n474), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n466), .B(new_n472), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(new_n470), .B2(G953), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(new_n468), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n461), .A2(new_n462), .A3(new_n455), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n454), .B(KEYINPUT8), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n321), .B1(new_n456), .B2(new_n458), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n234), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n461), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n479), .B1(new_n467), .B2(new_n468), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n477), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n477), .A2(new_n490), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(KEYINPUT88), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT84), .Z(new_n498));
  NAND2_X1  g312(.A1(G234), .A2(G237), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G952), .A3(new_n187), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT97), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT21), .B(G898), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n499), .A2(G902), .A3(G953), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n496), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(G104), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n211), .ZN(new_n512));
  NOR2_X1   g326(.A1(KEYINPUT89), .A2(G143), .ZN(new_n513));
  OAI211_X1 g327(.A(G214), .B(new_n343), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n343), .A2(G214), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n511), .B2(new_n211), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT18), .A2(G131), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n383), .B(new_n209), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n309), .B1(new_n514), .B2(new_n516), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n518), .B(new_n519), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n383), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n209), .C1(new_n383), .C2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n516), .A3(new_n309), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n387), .C1(new_n529), .C2(new_n520), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n510), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n309), .C1(new_n514), .C2(new_n516), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n421), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n532), .A3(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n520), .A2(KEYINPUT18), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n519), .A2(new_n518), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n531), .B1(new_n538), .B2(new_n510), .ZN(new_n539));
  NOR2_X1   g353(.A1(G475), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT20), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n520), .A2(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n420), .A3(new_n387), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n529), .A2(new_n520), .A3(KEYINPUT17), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n510), .B(new_n523), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n523), .A2(new_n530), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(new_n510), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n540), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n207), .B2(G143), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n211), .A2(KEYINPUT93), .A3(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n207), .A2(G143), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n246), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n246), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n556), .A2(new_n557), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G134), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT95), .A3(new_n558), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n318), .A2(G122), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n566));
  INV_X1    g380(.A(G122), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(G116), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n318), .A2(KEYINPUT92), .A3(G122), .ZN(new_n569));
  OAI221_X1 g383(.A(new_n565), .B1(KEYINPUT14), .B2(new_n198), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT14), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(G107), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n561), .A2(new_n564), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n556), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n554), .A2(KEYINPUT13), .A3(new_n555), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n557), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G134), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(G107), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n198), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n579), .A2(new_n580), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n298), .A2(new_n445), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n574), .A2(new_n585), .A3(new_n587), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT15), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G478), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n574), .A2(new_n585), .A3(new_n587), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n574), .B2(new_n585), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n592), .B(new_n289), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n593), .A3(G478), .ZN(new_n599));
  INV_X1    g413(.A(new_n546), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n535), .A2(new_n436), .A3(new_n543), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n510), .B1(new_n601), .B2(new_n523), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n289), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G475), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n551), .A2(new_n595), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n507), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n307), .A2(new_n382), .A3(new_n453), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n362), .B2(new_n289), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n362), .B2(new_n363), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n307), .A2(new_n453), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n497), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n477), .A2(new_n490), .ZN(new_n614));
  INV_X1    g428(.A(new_n491), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(new_n492), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n506), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n596), .B2(new_n597), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(KEYINPUT98), .B(new_n619), .C1(new_n596), .C2(new_n597), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n589), .A2(KEYINPUT33), .A3(new_n590), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n589), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n590), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n551), .A2(new_n604), .ZN(new_n632));
  INV_X1    g446(.A(G478), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n289), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n591), .B2(new_n633), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n618), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n612), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AOI22_X1  g454(.A1(new_n542), .A2(new_n550), .B1(G475), .B2(new_n603), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n599), .A2(new_n595), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n618), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n612), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n429), .A2(KEYINPUT36), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n418), .A2(new_n426), .A3(new_n648), .ZN(new_n649));
  OAI22_X1  g463(.A1(new_n435), .A2(new_n438), .B1(KEYINPUT36), .B2(new_n429), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n650), .A3(new_n450), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n440), .A2(new_n442), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n448), .A2(new_n447), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n449), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n307), .A2(new_n611), .A3(new_n606), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n504), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n501), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n641), .A2(new_n642), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n449), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT100), .B1(new_n449), .B2(new_n651), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n666), .B(new_n617), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n306), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n305), .B1(new_n296), .B2(new_n302), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n670), .B(new_n382), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n496), .B(KEYINPUT38), .Z(new_n675));
  NAND3_X1  g489(.A1(new_n632), .A2(new_n497), .A3(new_n642), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n675), .A2(new_n658), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n289), .B1(new_n374), .B2(new_n347), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n350), .B1(new_n339), .B2(new_n341), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n682), .B(G472), .C1(new_n678), .C2(new_n679), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n367), .A2(new_n381), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n664), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n307), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n677), .B(new_n685), .C1(new_n687), .C2(KEYINPUT40), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(KEYINPUT40), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n211), .ZN(G45));
  OAI21_X1  g504(.A(new_n617), .B1(new_n667), .B2(new_n668), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n631), .A2(new_n632), .A3(new_n635), .A4(new_n665), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n693), .B(new_n382), .C1(new_n671), .C2(new_n672), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n287), .A2(new_n289), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  INV_X1    g511(.A(new_n300), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n697), .A2(new_n290), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n382), .A2(new_n637), .A3(new_n453), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n382), .A2(new_n644), .A3(new_n453), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  INV_X1    g518(.A(new_n605), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n617), .B(new_n705), .C1(new_n667), .C2(new_n668), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n697), .A2(new_n290), .A3(new_n698), .A4(new_n506), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n708), .A2(KEYINPUT102), .A3(new_n382), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT102), .B1(new_n708), .B2(new_n382), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n316), .ZN(G21));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n610), .B(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n617), .A2(new_n715), .A3(new_n642), .A4(new_n632), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n477), .A2(new_n490), .A3(new_n491), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n491), .B1(new_n477), .B2(new_n490), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n497), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n632), .A2(new_n642), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT104), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n707), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n349), .B(new_n361), .C1(new_n347), .C2(new_n375), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n363), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n714), .A2(new_n722), .A3(new_n452), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT105), .B(G122), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G24));
  NAND2_X1  g541(.A1(new_n362), .A2(new_n289), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n713), .B1(new_n728), .B2(G472), .ZN(new_n729));
  AOI211_X1 g543(.A(KEYINPUT103), .B(new_n609), .C1(new_n362), .C2(new_n289), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n658), .B(new_n724), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n692), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n617), .A3(new_n699), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n492), .B(new_n497), .C1(new_n493), .C2(new_n495), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n291), .A2(new_n740), .A3(new_n293), .A4(G469), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n294), .A2(KEYINPUT106), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n290), .A2(new_n295), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n698), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT107), .A3(new_n698), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n382), .A3(new_n453), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n738), .B1(new_n748), .B2(new_n692), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(new_n745), .ZN(new_n750));
  INV_X1    g564(.A(new_n739), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n452), .ZN(new_n753));
  INV_X1    g567(.A(new_n381), .ZN(new_n754));
  INV_X1    g568(.A(new_n358), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n356), .A2(new_n341), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n347), .C1(new_n756), .C2(new_n351), .ZN(new_n757));
  INV_X1    g571(.A(new_n369), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n376), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n375), .B2(new_n377), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n609), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT32), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n364), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n753), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n752), .A2(new_n765), .A3(KEYINPUT42), .A4(new_n733), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n749), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  XOR2_X1   g582(.A(new_n666), .B(KEYINPUT108), .Z(new_n769));
  NOR2_X1   g583(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n246), .ZN(G36));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n611), .B1(new_n656), .B2(new_n657), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n631), .A2(new_n641), .A3(new_n635), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(KEYINPUT109), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT109), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n772), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n778), .A2(new_n779), .ZN(new_n783));
  INV_X1    g597(.A(new_n781), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT44), .A4(new_n774), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT45), .B1(new_n291), .B2(new_n293), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n288), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n291), .A2(KEYINPUT45), .A3(new_n293), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n295), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n290), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n698), .B(new_n686), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n739), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n782), .A2(new_n785), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  OAI21_X1  g610(.A(new_n698), .B1(new_n791), .B2(new_n792), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT47), .B(new_n698), .C1(new_n791), .C2(new_n792), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n382), .A2(new_n453), .A3(new_n692), .A4(new_n739), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(G140), .Z(G42));
  NAND2_X1  g618(.A1(new_n697), .A2(new_n290), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n452), .A2(new_n302), .A3(new_n498), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n806), .A2(new_n807), .A3(new_n775), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n685), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n675), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n776), .A2(new_n777), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n452), .B(new_n724), .C1(new_n729), .C2(new_n730), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n813), .A3(new_n501), .ZN(new_n814));
  INV_X1    g628(.A(new_n699), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n497), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n675), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT50), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(KEYINPUT50), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n815), .A2(new_n501), .A3(new_n739), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n823), .B2(new_n812), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(KEYINPUT116), .A3(new_n777), .A4(new_n776), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n822), .A2(new_n453), .A3(new_n810), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n632), .B1(new_n631), .B2(new_n635), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n826), .A2(new_n732), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n819), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n814), .A2(new_n751), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n697), .A2(new_n290), .A3(new_n301), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT114), .Z(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n801), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT51), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n826), .A2(new_n765), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT48), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n799), .A2(new_n800), .A3(new_n832), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n819), .A2(new_n840), .A3(new_n820), .A4(new_n829), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n814), .A2(new_n617), .A3(new_n699), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT117), .ZN(new_n843));
  INV_X1    g657(.A(G952), .ZN(new_n844));
  INV_X1    g658(.A(new_n636), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n844), .B(G953), .C1(new_n827), .C2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n837), .A2(new_n841), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n835), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n605), .B2(new_n664), .ZN(new_n850));
  INV_X1    g664(.A(new_n642), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT111), .A3(new_n641), .A4(new_n665), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n658), .A2(new_n850), .A3(new_n751), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n307), .A2(new_n853), .A3(new_n382), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n748), .B2(new_n769), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n746), .A2(new_n733), .A3(new_n747), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n731), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n767), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n507), .B1(new_n636), .B2(new_n643), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n307), .A2(new_n611), .A3(new_n453), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n607), .A2(new_n659), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT102), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n719), .B1(new_n656), .B2(new_n657), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n699), .A3(new_n506), .A4(new_n705), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n754), .A2(new_n761), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n863), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n708), .A2(KEYINPUT102), .A3(new_n382), .ZN(new_n869));
  INV_X1    g683(.A(new_n813), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n722), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n700), .A2(new_n703), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n862), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n859), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n716), .A2(new_n721), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n449), .A2(new_n651), .A3(new_n665), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n744), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n685), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n694), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n673), .A4(new_n736), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n673), .B1(new_n731), .B2(new_n734), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n694), .A2(new_n879), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n882), .B1(new_n881), .B2(new_n886), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n875), .B(KEYINPUT53), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n725), .B1(new_n709), .B2(new_n710), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n872), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n767), .A3(new_n862), .A4(new_n858), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  INV_X1    g708(.A(new_n673), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n731), .A2(new_n734), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(new_n897), .B2(new_n880), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n884), .A2(new_n885), .A3(new_n883), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n881), .A2(KEYINPUT112), .A3(new_n886), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n890), .B1(new_n902), .B2(KEYINPUT53), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n881), .A2(KEYINPUT112), .A3(new_n886), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT112), .B1(new_n881), .B2(new_n886), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n875), .B(KEYINPUT53), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT113), .B1(new_n898), .B2(new_n899), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n893), .B1(new_n909), .B2(new_n887), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n907), .B(new_n908), .C1(new_n910), .C2(KEYINPUT53), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n848), .A2(new_n904), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n844), .A2(new_n187), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n811), .B1(new_n915), .B2(new_n916), .ZN(G75));
  OAI21_X1  g731(.A(new_n907), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G210), .A3(G902), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n472), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT55), .Z(new_n924));
  AOI21_X1  g738(.A(KEYINPUT119), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n926));
  INV_X1    g740(.A(new_n924), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n926), .B(new_n927), .C1(new_n919), .C2(new_n920), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n187), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n918), .A2(G902), .A3(new_n494), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n924), .A2(KEYINPUT56), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n929), .A2(new_n937), .ZN(G51));
  NAND2_X1  g752(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n911), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n295), .B(KEYINPUT57), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n287), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n789), .B(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n918), .A2(G902), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n930), .B1(new_n943), .B2(new_n945), .ZN(G54));
  AND4_X1   g760(.A1(KEYINPUT58), .A2(new_n918), .A3(G475), .A4(G902), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n931), .B1(new_n947), .B2(new_n548), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n548), .B2(new_n947), .ZN(G60));
  INV_X1    g763(.A(new_n630), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n634), .B(KEYINPUT59), .Z(new_n951));
  AND3_X1   g765(.A1(new_n940), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n904), .A2(new_n911), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n950), .B1(new_n953), .B2(new_n951), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n954), .A3(new_n930), .ZN(G63));
  XOR2_X1   g769(.A(new_n444), .B(KEYINPUT60), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n918), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n431), .A2(new_n439), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n649), .A2(new_n650), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n931), .C1(new_n960), .C2(new_n957), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n503), .B2(new_n470), .ZN(new_n964));
  INV_X1    g778(.A(new_n874), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n922), .B1(G898), .B2(new_n187), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  OAI21_X1  g782(.A(new_n313), .B1(new_n338), .B2(KEYINPUT30), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT122), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n525), .B1(new_n383), .B2(new_n526), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n765), .A2(new_n876), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n793), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n803), .A2(new_n770), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n897), .A2(new_n694), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n976), .A2(new_n767), .A3(new_n795), .A4(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n972), .B(new_n973), .C1(new_n979), .C2(G953), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT62), .B1(new_n689), .B2(new_n977), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT123), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n739), .B1(new_n636), .B2(new_n643), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n382), .A3(new_n453), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n687), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n803), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n795), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n689), .A2(KEYINPUT62), .A3(new_n977), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(G953), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n980), .B1(new_n990), .B2(new_n972), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n980), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n991), .B(new_n994), .Z(G72));
  INV_X1    g809(.A(new_n679), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n339), .A2(new_n341), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(new_n347), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n903), .A2(new_n996), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT127), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n979), .B2(new_n874), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n930), .B1(new_n1005), .B2(new_n998), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n982), .A2(new_n989), .A3(new_n965), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1007), .A2(new_n1008), .A3(new_n1002), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n679), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1004), .A2(new_n1012), .ZN(G57));
endmodule


