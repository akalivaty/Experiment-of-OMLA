//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  XNOR2_X1  g000(.A(KEYINPUT85), .B(G36gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n203), .A2(KEYINPUT86), .A3(new_n205), .A4(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211));
  NAND2_X1  g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT84), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(KEYINPUT84), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(new_n205), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n220), .B1(G29gat), .B2(new_n202), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT86), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  INV_X1    g023(.A(new_n215), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT87), .B(KEYINPUT15), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n221), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT88), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n217), .A2(new_n222), .B1(new_n221), .B2(new_n227), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT88), .A3(new_n224), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT16), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G8gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT89), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n237), .B(new_n239), .C1(new_n236), .C2(new_n235), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(KEYINPUT89), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n232), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT17), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT90), .Z(new_n249));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n242), .B2(new_n243), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n242), .A2(new_n243), .A3(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n232), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(new_n249), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n247), .A2(KEYINPUT18), .A3(new_n249), .A4(new_n254), .ZN(new_n258));
  INV_X1    g057(.A(new_n253), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n245), .A3(new_n251), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n249), .B(KEYINPUT13), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT82), .B(G197gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT11), .B(G169gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n271), .A3(new_n258), .A4(new_n263), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(KEYINPUT22), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n277), .B1(new_n284), .B2(KEYINPUT29), .ZN(new_n285));
  XOR2_X1   g084(.A(G141gat), .B(G148gat), .Z(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT2), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G155gat), .B(G162gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n291), .A3(new_n289), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n277), .A3(new_n294), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n284), .ZN(new_n300));
  AND4_X1   g099(.A1(G228gat), .A2(new_n296), .A3(G233gat), .A4(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n296), .A2(new_n300), .B1(G228gat), .B2(G233gat), .ZN(new_n302));
  OAI21_X1  g101(.A(G22gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT78), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT31), .B(G50gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n301), .A2(G22gat), .A3(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n303), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n304), .A2(new_n309), .A3(new_n303), .A4(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n284), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(G169gat), .ZN(new_n318));
  INV_X1    g117(.A(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G183gat), .B(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n322), .B2(KEYINPUT24), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n328));
  INV_X1    g127(.A(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n323), .A2(new_n327), .A3(KEYINPUT25), .A4(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n332));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(new_n329), .ZN(new_n334));
  OAI221_X1 g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .C1(new_n321), .C2(new_n316), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n318), .A2(new_n319), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(KEYINPUT26), .B2(new_n329), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n338), .A2(new_n340), .B1(KEYINPUT28), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT27), .B(G183gat), .Z(new_n346));
  OAI21_X1  g145(.A(KEYINPUT67), .B1(new_n346), .B2(G190gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n348), .B1(G183gat), .B2(G190gat), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n331), .A2(new_n336), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n315), .B1(new_n350), .B2(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n331), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(G226gat), .A3(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n314), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n356), .A2(new_n284), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT30), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT0), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n295), .A2(KEYINPUT3), .ZN(new_n372));
  INV_X1    g171(.A(G113gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G120gat), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT69), .B(G120gat), .Z(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n373), .ZN(new_n376));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT1), .B1(new_n377), .B2(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n377), .ZN(new_n381));
  XNOR2_X1  g180(.A(G113gat), .B(G120gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT68), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n382), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n388), .A3(new_n297), .ZN(new_n389));
  INV_X1    g188(.A(new_n295), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n387), .A3(new_n380), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n388), .A2(new_n295), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n380), .A2(new_n387), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n390), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n396), .A2(new_n397), .B1(new_n402), .B2(KEYINPUT5), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n371), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(new_n397), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n371), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n413));
  INV_X1    g212(.A(new_n371), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n414), .A3(new_n410), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n406), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT6), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n367), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT74), .B1(new_n360), .B2(new_n361), .ZN(new_n420));
  INV_X1    g219(.A(new_n359), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT73), .B1(new_n351), .B2(new_n355), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n284), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n424));
  INV_X1    g223(.A(new_n361), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n365), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n360), .A2(new_n361), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(KEYINPUT75), .A3(KEYINPUT30), .A4(new_n364), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT30), .A4(new_n364), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n429), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n419), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT76), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n313), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n354), .A2(new_n400), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n350), .A2(new_n388), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(G227gat), .A4(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n442), .B(KEYINPUT32), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n442), .B2(KEYINPUT32), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n442), .A2(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT71), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n453), .A3(new_n450), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n448), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT34), .Z(new_n459));
  OAI21_X1  g258(.A(new_n439), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n449), .A2(new_n453), .A3(new_n450), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n453), .B1(new_n449), .B2(new_n450), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n447), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n459), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT72), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n455), .A2(new_n459), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT79), .B1(new_n438), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(KEYINPUT36), .B2(new_n467), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n437), .A2(new_n434), .A3(new_n419), .ZN(new_n476));
  INV_X1    g275(.A(new_n313), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n396), .A2(new_n397), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n401), .A2(new_n399), .A3(new_n393), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n371), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n417), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n484), .A2(KEYINPUT40), .A3(new_n371), .A4(new_n485), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n428), .A2(new_n364), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n427), .A3(new_n429), .A4(new_n433), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n477), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n416), .A2(new_n418), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n364), .B1(new_n428), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n314), .B1(new_n421), .B2(new_n422), .ZN(new_n499));
  INV_X1    g298(.A(new_n356), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n500), .B2(new_n284), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n366), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n420), .A2(KEYINPUT37), .A3(new_n426), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n498), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n496), .B(new_n503), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n495), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n473), .A2(new_n480), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n460), .A2(new_n313), .A3(new_n465), .A4(new_n466), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT35), .B1(new_n476), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n496), .A2(new_n477), .A3(KEYINPUT35), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n470), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n494), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT81), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n276), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT8), .ZN(new_n523));
  NAND2_X1  g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G85gat), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT97), .ZN(new_n535));
  AOI22_X1  g334(.A1(KEYINPUT8), .A2(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n536), .A2(new_n532), .A3(new_n526), .A4(new_n530), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(KEYINPUT97), .A3(new_n533), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT41), .ZN(new_n541));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n245), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n245), .B2(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n234), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT98), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n540), .B1(new_n232), .B2(new_n224), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n231), .B2(new_n233), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552));
  NOR4_X1   g351(.A1(new_n551), .A2(new_n552), .A3(new_n543), .A4(new_n547), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n546), .B2(new_n548), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT99), .B(new_n547), .C1(new_n551), .C2(new_n543), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(G162gat), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n233), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT88), .B1(new_n232), .B2(new_n224), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n545), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n543), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n548), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n552), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n546), .A2(KEYINPUT98), .A3(new_n548), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(new_n288), .A3(new_n556), .A4(new_n557), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n542), .A2(new_n541), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT96), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G134gat), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n559), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n559), .B2(new_n568), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  OR2_X1    g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  INV_X1    g379(.A(G57gat), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n580), .B(G64gat), .C1(new_n581), .C2(KEYINPUT93), .ZN(new_n582));
  INV_X1    g381(.A(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT92), .B1(new_n583), .B2(G57gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n583), .A3(G57gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT94), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n579), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT95), .Z(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n259), .B(new_n251), .C1(new_n592), .C2(new_n591), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n599), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n598), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n574), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n544), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n534), .A2(new_n537), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n579), .C1(new_n589), .C2(new_n590), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT10), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT10), .B(new_n579), .C1(new_n589), .C2(new_n590), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT100), .B1(new_n612), .B2(new_n544), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n540), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n606), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n607), .A2(new_n609), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n615), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n614), .B1(new_n540), .B2(new_n611), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n618), .A3(new_n609), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G120gat), .B(G148gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT101), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n617), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n605), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n521), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n496), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n236), .ZN(G1324gat));
  OAI21_X1  g442(.A(G8gat), .B1(new_n640), .B2(new_n517), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  NAND4_X1  g446(.A1(new_n521), .A2(new_n494), .A3(new_n639), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(G1325gat));
  INV_X1    g450(.A(new_n640), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n516), .A2(new_n518), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n472), .A2(G15gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT104), .Z(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n652), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n313), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NOR2_X1   g460(.A1(new_n604), .A2(new_n638), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n574), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n521), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n641), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT45), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n572), .A2(new_n573), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n511), .B2(new_n520), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n510), .A2(new_n475), .A3(new_n478), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n520), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n672), .B2(new_n668), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n273), .A2(new_n675), .A3(new_n274), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n273), .B2(new_n274), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(new_n679), .A3(new_n662), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n641), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT45), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n681), .A3(new_n682), .ZN(G1328gat));
  NOR3_X1   g482(.A1(new_n665), .A2(new_n202), .A3(new_n517), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n202), .B1(new_n680), .B2(new_n517), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(G1329gat));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n472), .A3(new_n679), .A4(new_n662), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G43gat), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n665), .A2(G43gat), .A3(new_n653), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(G1330gat));
  INV_X1    g496(.A(G50gat), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n670), .A2(new_n673), .A3(new_n678), .A4(new_n663), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n477), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n477), .A2(new_n698), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n665), .A2(new_n704), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n700), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n701), .B1(new_n700), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  INV_X1    g507(.A(new_n638), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n605), .A2(new_n709), .A3(new_n679), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n672), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n641), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n581), .ZN(G1332gat));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n494), .B(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  NOR3_X1   g520(.A1(new_n711), .A2(G71gat), .A3(new_n653), .ZN(new_n722));
  INV_X1    g521(.A(new_n711), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n472), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(G71gat), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n477), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g528(.A1(new_n511), .A2(new_n520), .ZN(new_n730));
  INV_X1    g529(.A(new_n669), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n673), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n679), .A2(new_n604), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n638), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n734), .A2(new_n641), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n574), .B1(new_n671), .B2(new_n520), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n735), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n738), .B2(new_n735), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n638), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n496), .A2(new_n527), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n737), .A2(new_n527), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n716), .A2(G92gat), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n638), .B(new_n745), .C1(new_n739), .C2(new_n740), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n734), .A2(new_n716), .A3(new_n736), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n744), .B(new_n746), .C1(new_n747), .C2(new_n528), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  INV_X1    g548(.A(new_n736), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n733), .A3(new_n494), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n749), .B(new_n744), .C1(new_n752), .C2(new_n746), .ZN(new_n753));
  NOR4_X1   g552(.A1(new_n670), .A2(new_n673), .A3(new_n517), .A4(new_n736), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n746), .B1(new_n754), .B2(new_n528), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT110), .B1(new_n755), .B2(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n748), .B1(new_n753), .B2(new_n756), .ZN(G1337gat));
  NOR3_X1   g556(.A1(new_n734), .A2(new_n475), .A3(new_n736), .ZN(new_n758));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n654), .A2(new_n759), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n758), .A2(new_n759), .B1(new_n741), .B2(new_n760), .ZN(G1338gat));
  INV_X1    g560(.A(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n477), .A2(new_n762), .A3(new_n638), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT111), .Z(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n739), .B2(new_n740), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n734), .A2(new_n313), .A3(new_n736), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n762), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n765), .C1(new_n766), .C2(new_n762), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n261), .A2(new_n262), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n249), .B1(new_n247), .B2(new_n254), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n269), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n638), .A2(new_n274), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n619), .A2(new_n779), .A3(new_n626), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n616), .A2(new_n618), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n635), .A3(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n633), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n633), .A4(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n637), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n678), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n574), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(new_n274), .A3(new_n777), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n572), .A2(new_n573), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n787), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n604), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(new_n795), .B1(new_n639), .B2(new_n678), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n796), .A2(new_n641), .A3(new_n512), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n716), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n373), .A3(new_n679), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n796), .A2(new_n477), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n800), .A2(new_n496), .A3(new_n654), .A4(new_n716), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n276), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n373), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT113), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n799), .B(new_n805), .C1(new_n373), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1340gat));
  INV_X1    g606(.A(new_n375), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n808), .A3(new_n638), .ZN(new_n809));
  OAI21_X1  g608(.A(G120gat), .B1(new_n801), .B2(new_n709), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n798), .A2(new_n812), .A3(new_n604), .ZN(new_n813));
  OAI21_X1  g612(.A(G127gat), .B1(new_n801), .B2(new_n795), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1342gat));
  NOR3_X1   g614(.A1(new_n574), .A2(G134gat), .A3(new_n494), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n797), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(KEYINPUT56), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n801), .B2(new_n574), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n818), .B2(new_n820), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(G1343gat));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n472), .A2(new_n715), .A3(new_n641), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n477), .A2(KEYINPUT57), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n783), .A2(new_n784), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n786), .A2(new_n637), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n785), .A2(new_n832), .A3(new_n637), .A4(new_n786), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n275), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n668), .B1(new_n834), .B2(new_n778), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n793), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT117), .B(new_n668), .C1(new_n834), .C2(new_n778), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n795), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n574), .A2(new_n604), .A3(new_n709), .A4(new_n678), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n828), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n788), .A2(new_n574), .B1(new_n791), .B2(new_n792), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n840), .B1(new_n843), .B2(new_n604), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(new_n477), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n679), .B(new_n827), .C1(new_n841), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G141gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n472), .A2(new_n313), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(new_n496), .A3(new_n716), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n276), .A2(G141gat), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n826), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n826), .B1(new_n849), .B2(new_n850), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n275), .B(new_n827), .C1(new_n841), .C2(new_n845), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(G141gat), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(G141gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n851), .B1(new_n846), .B2(G141gat), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n860), .B(new_n861), .C1(new_n826), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n863), .ZN(G1344gat));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n827), .B1(new_n841), .B2(new_n845), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(G148gat), .C1(new_n866), .C2(new_n709), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n844), .A2(new_n477), .A3(new_n842), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n639), .A2(new_n276), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n791), .A2(new_n792), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n795), .B1(new_n870), .B2(new_n835), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n313), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n638), .B1(new_n827), .B2(KEYINPUT119), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(KEYINPUT119), .B2(new_n827), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G148gat), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT120), .B1(new_n877), .B2(KEYINPUT59), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n879), .B(new_n865), .C1(new_n876), .C2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n867), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n849), .A2(G148gat), .A3(new_n709), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n866), .B2(new_n795), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n604), .A2(new_n287), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n849), .B2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n866), .B2(new_n574), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n844), .A2(new_n496), .A3(new_n848), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n668), .A2(new_n288), .A3(new_n517), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n517), .A2(new_n496), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n653), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n800), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n318), .A3(new_n276), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n844), .A2(new_n641), .A3(new_n715), .ZN(new_n896));
  INV_X1    g695(.A(new_n512), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n679), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n895), .B1(new_n318), .B2(new_n898), .ZN(G1348gat));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n319), .B1(new_n900), .B2(new_n709), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT122), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n894), .A2(new_n319), .A3(new_n709), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1349gat));
  OAI21_X1  g703(.A(KEYINPUT124), .B1(new_n894), .B2(new_n795), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n800), .A2(new_n906), .A3(new_n604), .A4(new_n893), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(G183gat), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n795), .A2(new_n346), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n897), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n897), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n894), .B2(new_n574), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n668), .A2(new_n343), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n921), .A2(new_n922), .B1(new_n900), .B2(new_n923), .ZN(G1351gat));
  AND2_X1   g723(.A1(new_n896), .A2(new_n848), .ZN(new_n925));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n679), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n892), .A2(new_n472), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n873), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n275), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  AOI21_X1  g731(.A(G204gat), .B1(new_n932), .B2(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n638), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G204gat), .B1(new_n928), .B2(new_n709), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n925), .A2(new_n279), .A3(new_n604), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n873), .A2(new_n604), .A3(new_n927), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n873), .A2(new_n944), .A3(new_n604), .A4(new_n927), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(G211gat), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT63), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n943), .A2(new_n948), .A3(G211gat), .A4(new_n945), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n947), .A3(new_n949), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n928), .B2(new_n574), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n280), .A3(new_n668), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


