//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  OR3_X1    g0021(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n222));
  OAI21_X1  g0022(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n221), .B(new_n226), .C1(new_n229), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n209), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT67), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(G223), .A3(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n255), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G77), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  INV_X1    g0079(.A(G1), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n252), .B1(new_n270), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(KEYINPUT68), .B(new_n284), .C1(new_n268), .C2(new_n269), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G179), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n228), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G20), .B2(new_n203), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(new_n227), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n280), .A2(G13), .A3(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n227), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n280), .A2(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(G50), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G50), .B2(new_n301), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n286), .A2(new_n287), .A3(G169), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n290), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(G190), .B1(new_n286), .B2(new_n287), .ZN(new_n313));
  XOR2_X1   g0113(.A(new_n308), .B(KEYINPUT9), .Z(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n286), .A2(new_n287), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n313), .B(new_n314), .C1(new_n316), .C2(KEYINPUT72), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n288), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT10), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n314), .A2(new_n313), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n318), .B1(new_n288), .B2(new_n315), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n312), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n283), .A2(G1698), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G223), .B2(G1698), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n253), .A2(new_n254), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n257), .B2(new_n211), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n269), .B1(new_n274), .B2(new_n277), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT79), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n282), .B2(new_n216), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n279), .A2(KEYINPUT79), .A3(G232), .A4(new_n281), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n315), .B1(new_n331), .B2(new_n335), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n215), .A2(new_n209), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n341), .B2(new_n201), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n294), .A2(G159), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n258), .A2(new_n260), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n349), .B2(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n299), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(G20), .B1(new_n255), .B2(new_n261), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n352), .B2(KEYINPUT7), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n344), .B1(new_n353), .B2(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(KEYINPUT16), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n291), .B1(new_n280), .B2(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n304), .B1(new_n302), .B2(new_n291), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n340), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT17), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n340), .A2(new_n355), .A3(KEYINPUT17), .A4(new_n357), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G244), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n266), .A2(G107), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n278), .B1(new_n363), .B2(new_n282), .C1(new_n367), .C2(new_n279), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n304), .A2(G77), .A3(new_n305), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT70), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n304), .A2(new_n373), .A3(G77), .A4(new_n305), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n372), .A2(new_n374), .B1(new_n375), .B2(new_n302), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n291), .A2(new_n295), .B1(new_n228), .B2(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n377), .A2(new_n378), .B1(new_n292), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n303), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n370), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n368), .A2(G179), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n353), .A2(G68), .ZN(new_n387));
  INV_X1    g0187(.A(new_n344), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT16), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n346), .A2(new_n345), .A3(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n329), .B2(new_n228), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n388), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n303), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n357), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n336), .A2(G169), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n331), .A2(new_n335), .A3(G179), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT18), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n396), .A2(KEYINPUT80), .A3(KEYINPUT18), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n399), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n383), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n368), .A2(G200), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n337), .C2(new_n368), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n362), .A2(new_n386), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n278), .B1(new_n282), .B2(new_n210), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n255), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n255), .A2(new_n261), .A3(G226), .A4(new_n263), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n269), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n418), .A2(KEYINPUT74), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT74), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n269), .ZN(new_n423));
  INV_X1    g0223(.A(new_n413), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n418), .B2(new_n419), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n294), .A2(G50), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n432), .B(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n292), .A2(new_n375), .B1(new_n228), .B2(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n303), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT11), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT11), .B(new_n303), .C1(new_n434), .C2(new_n435), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT12), .B1(new_n301), .B2(G68), .ZN(new_n440));
  OR3_X1    g0240(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n209), .B1(new_n280), .B2(G20), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n440), .A2(new_n441), .B1(new_n304), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n418), .A2(new_n419), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n431), .B(new_n446), .C1(new_n315), .C2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n422), .A2(G179), .A3(new_n429), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n422), .A2(new_n429), .A3(KEYINPUT77), .A4(G179), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT14), .B1(new_n449), .B2(new_n369), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT14), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(G169), .C1(new_n447), .C2(new_n448), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT78), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n446), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n446), .A2(new_n462), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n326), .A2(new_n412), .A3(new_n450), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT4), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n363), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n255), .A2(new_n261), .A3(new_n263), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n255), .A2(new_n261), .A3(G250), .A4(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(new_n263), .C1(new_n253), .C2(new_n254), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n475), .A2(new_n469), .B1(G33), .B2(G283), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n269), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n276), .A2(G1), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n269), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n274), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(new_n486), .A3(new_n289), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n262), .A2(KEYINPUT81), .A3(new_n263), .A4(new_n470), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n491), .A2(new_n473), .A3(new_n474), .A4(new_n476), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n269), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n489), .A2(new_n369), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n490), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n353), .A2(G107), .ZN(new_n499));
  INV_X1    g0299(.A(G107), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  XOR2_X1   g0301(.A(G97), .B(G107), .Z(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n303), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n301), .A2(G97), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n280), .A2(G33), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n299), .A2(new_n301), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n495), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n489), .A2(G200), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n487), .B1(new_n492), .B2(new_n269), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n513), .A2(new_n506), .A3(new_n515), .A4(new_n510), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n228), .B1(new_n416), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n211), .A2(new_n217), .A3(new_n500), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n228), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n292), .B2(new_n217), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n303), .ZN(new_n524));
  INV_X1    g0324(.A(new_n379), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n509), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n379), .A2(new_n302), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n363), .A2(G1698), .ZN(new_n529));
  OAI221_X1 g0329(.A(new_n529), .B1(G238), .B2(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n279), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n274), .A2(new_n480), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n212), .B1(new_n280), .B2(G45), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n279), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n369), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n274), .A2(new_n480), .B1(new_n279), .B2(new_n534), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G238), .A2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n363), .B2(G1698), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n346), .B1(G33), .B2(G116), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n289), .B(new_n538), .C1(new_n541), .C2(new_n279), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n528), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(G200), .B1(new_n532), .B2(new_n536), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n523), .A2(new_n303), .B1(new_n302), .B2(new_n379), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n509), .A2(G87), .ZN(new_n546));
  OAI211_X1 g0346(.A(G190), .B(new_n538), .C1(new_n541), .C2(new_n279), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT83), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n543), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n512), .A2(new_n516), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n304), .A2(new_n508), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n500), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT25), .B1(new_n302), .B2(new_n500), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n555), .A2(new_n500), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n211), .A2(KEYINPUT22), .A3(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n255), .A2(new_n261), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n228), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n531), .B2(G20), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n228), .A2(KEYINPUT86), .A3(G33), .A4(G116), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n500), .A3(G20), .ZN(new_n572));
  NAND2_X1  g0372(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n565), .A2(new_n575), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT88), .B1(new_n581), .B2(new_n303), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n565), .A2(new_n575), .A3(new_n577), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n565), .B2(new_n575), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT88), .B(new_n303), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n560), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n484), .A2(G264), .A3(new_n279), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G250), .A2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n218), .B2(G1698), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n346), .B1(G33), .B2(G294), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n486), .B(new_n588), .C1(new_n279), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n289), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT89), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT89), .B1(new_n592), .B2(G169), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n303), .B1(new_n583), .B2(new_n584), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT88), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n559), .B1(new_n601), .B2(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(new_n315), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G190), .B2(new_n592), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n482), .A2(G270), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n486), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n266), .A2(G303), .ZN(new_n610));
  AND2_X1   g0410(.A1(G264), .A2(G1698), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n346), .A2(KEYINPUT84), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n263), .C1(new_n253), .C2(new_n254), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n253), .B2(new_n254), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n610), .A2(new_n612), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n609), .B1(new_n617), .B2(new_n269), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n302), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n555), .B2(new_n619), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n298), .A2(new_n227), .B1(G20), .B2(new_n619), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(G33), .B2(G283), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(G33), .B2(new_n217), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n622), .A2(new_n624), .A3(KEYINPUT20), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT20), .B1(new_n622), .B2(new_n624), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G169), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n607), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n616), .A2(new_n612), .A3(new_n613), .ZN(new_n630));
  INV_X1    g0430(.A(G303), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n255), .B2(new_n261), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n269), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n482), .A2(G270), .B1(new_n485), .B2(new_n274), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI221_X1 g0435(.A(new_n620), .B1(new_n555), .B2(new_n619), .C1(new_n625), .C2(new_n626), .ZN(new_n636));
  INV_X1    g0436(.A(new_n607), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(G169), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n618), .A2(G179), .A3(new_n636), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n635), .A2(new_n337), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n315), .B1(new_n633), .B2(new_n634), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n468), .A2(new_n554), .A3(new_n606), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n467), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n446), .B1(new_n315), .B2(new_n449), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n430), .B2(G190), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n386), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n362), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n396), .A2(KEYINPUT18), .A3(new_n399), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT18), .B1(new_n396), .B2(new_n399), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n320), .A2(new_n325), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n312), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n468), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n553), .A2(new_n498), .A3(new_n495), .A4(new_n511), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(new_n662));
  INV_X1    g0462(.A(new_n597), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n602), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n549), .B1(new_n602), .B2(new_n604), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n512), .A2(new_n516), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n543), .B(new_n661), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n489), .A2(new_n369), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n493), .A2(new_n494), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n498), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT90), .ZN(new_n672));
  INV_X1    g0472(.A(new_n549), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n495), .A2(new_n674), .A3(new_n498), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n511), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n659), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n658), .A2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n280), .A2(new_n228), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n636), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n644), .A2(new_n687), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT92), .B1(new_n690), .B2(new_n693), .ZN(new_n697));
  INV_X1    g0497(.A(new_n686), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n602), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n606), .A2(new_n699), .B1(new_n598), .B2(new_n698), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n696), .A2(new_n697), .A3(G330), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n640), .A2(new_n698), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n598), .A3(new_n605), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n598), .A2(new_n686), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n224), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n519), .A2(G116), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n710), .A2(new_n280), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n232), .B2(new_n710), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n698), .C1(new_n668), .C2(new_n677), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n512), .A2(new_n516), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n664), .A3(new_n665), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n543), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(KEYINPUT26), .B2(new_n676), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(KEYINPUT94), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n724), .B(new_n721), .C1(KEYINPUT26), .C2(new_n676), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n698), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n718), .B1(new_n726), .B2(KEYINPUT29), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n588), .B1(new_n591), .B2(new_n279), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n538), .B1(new_n541), .B2(new_n279), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(G179), .A3(new_n633), .A4(new_n634), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n728), .B1(new_n489), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n592), .A2(new_n289), .A3(new_n730), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n489), .A2(new_n635), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n633), .A2(G179), .A3(new_n634), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n532), .A2(new_n536), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n591), .A2(new_n279), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n588), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n733), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n686), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n598), .A2(new_n644), .A3(new_n605), .A4(new_n698), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n554), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n686), .A2(KEYINPUT31), .ZN(new_n748));
  INV_X1    g0548(.A(new_n741), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n733), .A2(new_n735), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n750), .B2(KEYINPUT93), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n733), .A2(new_n752), .A3(new_n735), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n748), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n727), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n715), .B1(new_n756), .B2(G1), .ZN(G364));
  INV_X1    g0557(.A(G13), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n280), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n710), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n262), .A2(G355), .A3(new_n224), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n709), .A2(new_n346), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n231), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n250), .A2(new_n276), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n764), .B1(G116), .B2(new_n224), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n227), .B1(G20), .B2(new_n369), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n763), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n228), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G159), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT32), .Z(new_n782));
  NAND3_X1  g0582(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n228), .B1(new_n778), .B2(G190), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n782), .B1(new_n209), .B2(new_n785), .C1(new_n217), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n777), .A2(new_n289), .A3(G200), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n500), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n228), .A2(new_n337), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n289), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n211), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n787), .A2(new_n266), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n289), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n777), .A2(new_n797), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G58), .A2(new_n799), .B1(new_n801), .B2(G77), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n783), .A2(new_n337), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n202), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT96), .Z(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n800), .A2(new_n807), .B1(new_n786), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G326), .B2(new_n803), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT98), .Z(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n262), .B1(new_n784), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n780), .A2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(new_n794), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G303), .B1(new_n799), .B2(G322), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n791), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G283), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n796), .A2(new_n806), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n774), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n776), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n696), .A2(new_n697), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n773), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n696), .A2(new_n697), .A3(G330), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n763), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G330), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n824), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n678), .A2(new_n698), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n384), .A2(new_n385), .A3(new_n686), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n383), .A2(new_n686), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n411), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n386), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n698), .B(new_n836), .C1(new_n668), .C2(new_n677), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n762), .B1(new_n840), .B2(new_n755), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n755), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n774), .A2(new_n769), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT99), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n763), .B1(new_n845), .B2(new_n375), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n818), .A2(G87), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n815), .A2(G107), .B1(new_n799), .B2(G294), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n801), .A2(G116), .B1(new_n780), .B2(G311), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n266), .B1(new_n217), .B2(new_n786), .ZN(new_n851));
  INV_X1    g0651(.A(G283), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n785), .A2(new_n852), .B1(new_n804), .B2(new_n631), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT100), .Z(new_n855));
  NAND2_X1  g0655(.A1(new_n818), .A2(G68), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n202), .B2(new_n794), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  AOI22_X1  g0658(.A1(G143), .A2(new_n799), .B1(new_n801), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n804), .B2(new_n860), .C1(new_n293), .C2(new_n785), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n329), .B1(new_n780), .B2(G132), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n215), .B2(new_n786), .ZN(new_n866));
  OR3_X1    g0666(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n855), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n774), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n846), .B1(new_n770), .B2(new_n836), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n842), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(G384));
  NOR2_X1   g0674(.A1(new_n759), .A2(new_n280), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n466), .B(new_n686), .C1(new_n461), .C2(new_n649), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n463), .A2(new_n464), .A3(new_n686), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n459), .B1(new_n453), .B2(new_n454), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n450), .B(new_n877), .C1(new_n878), .C2(new_n465), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n745), .B(new_n881), .C1(new_n746), .C2(new_n554), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n880), .A2(new_n836), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(new_n684), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n396), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n404), .A2(new_n887), .A3(new_n358), .A4(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n404), .A2(new_n887), .A3(new_n358), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n360), .B(new_n361), .C1(new_n652), .C2(new_n653), .ZN(new_n894));
  INV_X1    g0694(.A(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n890), .A2(new_n892), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n358), .ZN(new_n900));
  INV_X1    g0700(.A(new_n399), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n351), .B1(KEYINPUT16), .B2(new_n350), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n684), .B1(new_n902), .B2(new_n357), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n889), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n407), .A2(new_n362), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n357), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n886), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT38), .B(new_n905), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n884), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n407), .B2(new_n362), .ZN(new_n911));
  INV_X1    g0711(.A(new_n905), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n885), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n914), .A2(new_n836), .A3(new_n880), .A4(new_n882), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n883), .A2(new_n910), .B1(new_n915), .B2(new_n884), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n659), .B2(new_n882), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n828), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n659), .A3(new_n882), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT105), .Z(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n833), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n839), .A2(new_n923), .B1(new_n879), .B2(new_n876), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n914), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n654), .A2(new_n684), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT39), .B1(new_n899), .B2(new_n909), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n467), .A2(new_n686), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n658), .B1(new_n727), .B2(new_n468), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n875), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n922), .B2(new_n935), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n938), .A2(G116), .A3(new_n229), .A4(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(G77), .B1(new_n215), .B2(new_n209), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n246), .B1(new_n231), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(G1), .A3(new_n758), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n942), .A3(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n775), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n709), .B2(new_n525), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n765), .A2(new_n241), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n763), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n543), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n698), .B1(new_n545), .B2(new_n546), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n549), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n794), .A2(new_n619), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(KEYINPUT46), .B1(new_n500), .B2(new_n786), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G311), .B2(new_n803), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n800), .A2(new_n852), .B1(new_n779), .B2(new_n958), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n346), .B(new_n959), .C1(G303), .C2(new_n799), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n818), .A2(G97), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n955), .A2(KEYINPUT46), .B1(new_n784), .B2(G294), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n818), .A2(G77), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n266), .B1(new_n784), .B2(G159), .ZN(new_n965));
  INV_X1    g0765(.A(new_n786), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n966), .A2(G68), .B1(G143), .B2(new_n803), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n794), .A2(new_n215), .B1(new_n800), .B2(new_n202), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n798), .A2(new_n293), .B1(new_n779), .B2(new_n860), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n965), .A3(new_n967), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n963), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT107), .Z(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n950), .B1(new_n772), .B2(new_n954), .C1(new_n974), .C2(new_n821), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n511), .A2(new_n686), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n719), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n672), .A2(new_n511), .A3(new_n675), .A4(new_n686), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n701), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n977), .A2(new_n978), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n705), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n598), .B1(new_n977), .B2(new_n978), .ZN(new_n988));
  INV_X1    g0788(.A(new_n512), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n698), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT106), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n987), .B2(new_n990), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n983), .B(new_n984), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT43), .A4(new_n954), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n981), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n984), .B1(new_n994), .B2(new_n995), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n982), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n980), .A3(new_n996), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n704), .B1(new_n700), .B2(new_n703), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n825), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n704), .B1(new_n598), .B2(new_n686), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT44), .B1(new_n979), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n707), .A2(new_n985), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n707), .A2(new_n985), .A3(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT45), .B1(new_n707), .B2(new_n985), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1007), .A2(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n701), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n979), .B2(new_n1006), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n707), .A2(new_n985), .A3(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n1006), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1008), .B1(new_n707), .B2(new_n985), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1021), .A3(new_n701), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n756), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n710), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n761), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n975), .B1(new_n1003), .B2(new_n1027), .ZN(G387));
  XOR2_X1   g0828(.A(new_n825), .B(new_n1004), .Z(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n727), .A3(new_n755), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n727), .A2(new_n755), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1032), .A3(new_n710), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n765), .B1(new_n238), .B2(new_n276), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n262), .A2(new_n224), .A3(new_n712), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n291), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT50), .B1(new_n291), .B2(G50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1037), .A2(new_n711), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(new_n500), .B2(new_n709), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n762), .B1(new_n1041), .B2(new_n947), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G317), .A2(new_n799), .B1(new_n801), .B2(G303), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT108), .B(G322), .Z(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n804), .B2(new_n1044), .C1(new_n807), .C2(new_n785), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n815), .A2(G294), .B1(new_n966), .B2(G283), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n818), .A2(G116), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n346), .B1(new_n780), .B2(G326), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n346), .B1(new_n779), .B2(new_n293), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n525), .B2(new_n966), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n291), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1059), .A2(new_n784), .B1(G159), .B2(new_n803), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n794), .A2(new_n375), .B1(new_n798), .B2(new_n202), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G68), .B2(new_n801), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n961), .A2(new_n1058), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n821), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n700), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1042), .B(new_n1064), .C1(new_n1065), .C2(new_n773), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1029), .B2(new_n761), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1033), .A2(new_n1067), .ZN(G393));
  AND3_X1   g0868(.A1(new_n1018), .A2(new_n701), .A3(new_n1021), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n701), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n761), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n775), .B1(new_n217), .B2(new_n224), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n245), .A2(new_n709), .A3(new_n346), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n762), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n799), .A2(G311), .B1(G317), .B2(new_n803), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n266), .B1(new_n619), .B2(new_n786), .C1(new_n631), .C2(new_n785), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n801), .A2(G294), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n852), .B2(new_n794), .C1(new_n779), .C2(new_n1044), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1077), .A2(new_n792), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT109), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n799), .A2(G159), .B1(G150), .B2(new_n803), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n346), .B1(new_n800), .B2(new_n291), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n794), .A2(new_n209), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G143), .C2(new_n780), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n786), .A2(new_n375), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n784), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n847), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1082), .A2(KEYINPUT109), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1083), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1075), .B1(new_n1093), .B2(new_n774), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n985), .B2(new_n772), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1072), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n710), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n1071), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1030), .A2(new_n1023), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  OAI22_X1  g0902(.A1(new_n928), .A2(new_n929), .B1(new_n924), .B2(new_n931), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n880), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n835), .A2(new_n386), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n698), .B(new_n1105), .C1(new_n723), .C2(new_n725), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n923), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n899), .A2(new_n909), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n467), .B2(new_n686), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n882), .A2(G330), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n880), .A2(new_n1112), .A3(new_n836), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n836), .C1(new_n747), .C2(new_n754), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n880), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1103), .B(new_n1118), .C1(new_n1107), .C2(new_n1109), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1106), .A2(new_n923), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1111), .A2(new_n837), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1118), .B1(new_n880), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT111), .B1(new_n1117), .B2(new_n880), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT111), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1116), .A2(new_n1126), .A3(new_n879), .A4(new_n876), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1113), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n839), .A2(new_n923), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT112), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT112), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1124), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n659), .A2(KEYINPUT110), .A3(new_n1112), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT110), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n468), .B2(new_n1111), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n658), .C1(new_n727), .C2(new_n468), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1120), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1124), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1128), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1132), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1139), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1119), .A3(new_n1115), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1146), .A3(new_n710), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1120), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n769), .B1(new_n928), .B2(new_n929), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n762), .B1(new_n844), .B2(new_n1059), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n785), .A2(new_n860), .B1(new_n804), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n266), .B(new_n1152), .C1(G159), .C2(new_n966), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n818), .A2(G50), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n799), .A2(G132), .B1(new_n801), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n779), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n794), .A2(new_n293), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1153), .A2(new_n1154), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n856), .B1(new_n808), .B2(new_n779), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT115), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT115), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n798), .A2(new_n619), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n262), .A2(new_n795), .A3(new_n1167), .A4(new_n1089), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n785), .A2(new_n500), .B1(new_n800), .B2(new_n217), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT113), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1170), .A2(new_n1171), .B1(new_n852), .B2(new_n804), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT114), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1163), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1150), .B1(new_n1175), .B2(new_n774), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1148), .A2(new_n761), .B1(new_n1149), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1147), .A2(new_n1177), .ZN(G378));
  NOR2_X1   g0978(.A1(new_n346), .A2(G41), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G50), .B(new_n1179), .C1(new_n257), .C2(new_n275), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n780), .A2(G283), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n379), .B2(new_n800), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1179), .B1(new_n794), .B2(new_n375), .C1(new_n217), .C2(new_n785), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G107), .C2(new_n799), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n804), .A2(new_n619), .B1(new_n786), .B2(new_n209), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT116), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n818), .A2(G58), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT117), .Z(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1180), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n794), .A2(new_n1155), .B1(new_n798), .B2(new_n1151), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n966), .A2(G150), .B1(G132), .B2(new_n784), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1158), .B2(new_n804), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G137), .C2(new_n801), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT59), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT118), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT118), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n818), .A2(G159), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1191), .B1(new_n1190), .B2(new_n1189), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n774), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT119), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n763), .B1(new_n202), .B2(new_n843), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n308), .A2(new_n684), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n326), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n326), .A2(new_n1210), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n326), .A2(new_n1210), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1211), .A3(new_n1207), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1206), .B1(new_n769), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n916), .B2(G330), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n915), .A2(new_n884), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n883), .A2(new_n910), .ZN(new_n1222));
  AND4_X1   g1022(.A1(G330), .A2(new_n1217), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n933), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1221), .A3(G330), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1218), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n916), .A2(G330), .A3(new_n1217), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n932), .A4(new_n927), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1219), .B1(new_n1229), .B2(new_n761), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1145), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(KEYINPUT57), .A3(new_n1229), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n710), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1229), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1230), .B1(new_n1233), .B2(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1141), .B(new_n1139), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1026), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1104), .A2(new_n769), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n798), .A2(new_n860), .B1(new_n800), .B2(new_n293), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G159), .B2(new_n815), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n346), .B1(new_n779), .B2(new_n1151), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G50), .B2(new_n966), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1156), .A2(new_n784), .B1(G132), .B2(new_n803), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1187), .A2(new_n1241), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n262), .B1(new_n525), .B2(new_n966), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n794), .A2(new_n217), .B1(new_n779), .B2(new_n631), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n798), .A2(new_n852), .B1(new_n800), .B2(new_n500), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n784), .A2(G116), .B1(new_n803), .B2(G294), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n964), .A2(new_n1246), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n821), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n763), .B(new_n1252), .C1(new_n209), .C2(new_n845), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1144), .A2(new_n761), .B1(new_n1239), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1238), .A2(new_n1254), .ZN(G381));
  OR2_X1    g1055(.A1(G375), .A2(G378), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1031), .B1(new_n1071), .B2(new_n1029), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n760), .B1(new_n1257), .B2(new_n1025), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1002), .A3(new_n999), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n975), .A3(new_n1101), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1033), .A2(new_n830), .A3(new_n1067), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n873), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT120), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G381), .A2(new_n1256), .A3(new_n1260), .A4(new_n1264), .ZN(G407));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  OAI211_X1 g1066(.A(G378), .B(new_n1230), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1267));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1231), .A2(new_n1026), .A3(new_n1229), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1230), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1097), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT60), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1237), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT121), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1273), .A2(new_n1277), .A3(new_n1275), .A4(KEYINPUT121), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1254), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n873), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n685), .A2(G213), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(G384), .A3(new_n1254), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1272), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n685), .A2(G213), .A3(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1284), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1272), .A2(new_n1285), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1282), .B2(new_n1254), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1254), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n873), .B(new_n1294), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1292), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1290), .A2(new_n1291), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1267), .A2(new_n1271), .B1(G213), .B2(new_n685), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1288), .A2(new_n1297), .A3(new_n1298), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT122), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n830), .B1(new_n1033), .B2(new_n1067), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1262), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(G387), .A2(G390), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1101), .B1(new_n1259), .B2(new_n975), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1304), .B(new_n1306), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(G390), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT122), .B1(new_n1262), .B2(new_n1305), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1305), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1304), .A3(new_n1261), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .A4(new_n1260), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT124), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1309), .A2(KEYINPUT124), .A3(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1303), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1309), .A2(new_n1298), .A3(new_n1314), .ZN(new_n1322));
  XOR2_X1   g1122(.A(new_n1322), .B(KEYINPUT123), .Z(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1287), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1299), .A2(new_n1300), .A3(KEYINPUT63), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1323), .A2(new_n1325), .A3(new_n1297), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1321), .A2(new_n1327), .ZN(G405));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1268), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1267), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1300), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1334), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1331), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1329), .B(new_n1320), .C1(new_n1335), .C2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1320), .A2(new_n1329), .ZN(new_n1340));
  AOI22_X1  g1140(.A1(new_n1319), .A2(KEYINPUT126), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1293), .A2(new_n1295), .A3(KEYINPUT125), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1337), .B1(new_n1336), .B2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1341), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(G402));
endmodule


