

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X2 U325 ( .A(n434), .B(KEYINPUT64), .Z(n570) );
  NOR2_X2 U326 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n453), .B(n452), .ZN(n528) );
  NOR2_X1 U328 ( .A1(n454), .A2(n528), .ZN(n566) );
  XNOR2_X1 U329 ( .A(n477), .B(KEYINPUT38), .ZN(n500) );
  XOR2_X1 U330 ( .A(n452), .B(n408), .Z(n518) );
  XOR2_X1 U331 ( .A(G190GAT), .B(KEYINPUT80), .Z(n401) );
  XNOR2_X1 U332 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U333 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U334 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U335 ( .A(n399), .B(n398), .ZN(n405) );
  XNOR2_X1 U336 ( .A(n558), .B(KEYINPUT36), .ZN(n584) );
  INV_X1 U337 ( .A(n380), .ZN(n381) );
  INV_X1 U338 ( .A(n558), .ZN(n565) );
  XNOR2_X1 U339 ( .A(n382), .B(n381), .ZN(n558) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n478), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT21), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(G197GAT), .B(n295), .Z(n399) );
  XOR2_X1 U348 ( .A(KEYINPUT76), .B(G162GAT), .Z(n373) );
  XOR2_X1 U349 ( .A(G78GAT), .B(G148GAT), .Z(n297) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n342) );
  XOR2_X1 U352 ( .A(n373), .B(n342), .Z(n299) );
  NAND2_X1 U353 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n399), .B(n300), .ZN(n312) );
  XOR2_X1 U356 ( .A(G204GAT), .B(KEYINPUT92), .Z(n302) );
  XNOR2_X1 U357 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U359 ( .A(n303), .B(KEYINPUT91), .Z(n305) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G22GAT), .Z(n324) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(n324), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n306), .B(KEYINPUT22), .Z(n310) );
  XOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT3), .Z(n308) );
  XNOR2_X1 U365 ( .A(KEYINPUT2), .B(KEYINPUT90), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n420) );
  XNOR2_X1 U367 ( .A(n420), .B(KEYINPUT23), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n470) );
  XOR2_X1 U370 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n386) );
  XNOR2_X1 U371 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n313), .B(G29GAT), .ZN(n314) );
  XOR2_X1 U373 ( .A(n314), .B(KEYINPUT8), .Z(n316) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G50GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n379) );
  XNOR2_X1 U376 ( .A(G15GAT), .B(G1GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n317), .B(KEYINPUT67), .ZN(n346) );
  XOR2_X1 U378 ( .A(n346), .B(KEYINPUT29), .Z(n319) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U381 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n321) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(G197GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U384 ( .A(n323), .B(n322), .Z(n326) );
  XOR2_X1 U385 ( .A(G169GAT), .B(G8GAT), .Z(n400) );
  XNOR2_X1 U386 ( .A(n324), .B(n400), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U388 ( .A(n379), .B(n327), .Z(n546) );
  INV_X1 U389 ( .A(n546), .ZN(n571) );
  XOR2_X1 U390 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n329) );
  XNOR2_X1 U391 ( .A(KEYINPUT75), .B(KEYINPUT69), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U393 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n331) );
  XOR2_X1 U394 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT13), .Z(n347) );
  XNOR2_X1 U396 ( .A(n443), .B(n347), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U401 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n337) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U404 ( .A(G85GAT), .B(n338), .Z(n380) );
  XOR2_X1 U405 ( .A(n339), .B(n380), .Z(n344) );
  XOR2_X1 U406 ( .A(G64GAT), .B(KEYINPUT74), .Z(n341) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n397) );
  XNOR2_X1 U409 ( .A(n342), .B(n397), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n344), .B(n343), .ZN(n577) );
  XOR2_X1 U411 ( .A(KEYINPUT41), .B(n577), .Z(n455) );
  AND2_X1 U412 ( .A1(n571), .A2(n455), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n345), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U414 ( .A(n347), .B(n346), .Z(n349) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n365) );
  XOR2_X1 U417 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n351) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n363) );
  XOR2_X1 U420 ( .A(G155GAT), .B(G71GAT), .Z(n353) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(G127GAT), .ZN(n352) );
  XNOR2_X1 U422 ( .A(n353), .B(n352), .ZN(n361) );
  XOR2_X1 U423 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n355) );
  XNOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U426 ( .A(G64GAT), .B(G78GAT), .Z(n357) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U429 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U431 ( .A(n363), .B(n362), .Z(n364) );
  XOR2_X1 U432 ( .A(n365), .B(n364), .Z(n555) );
  INV_X1 U433 ( .A(n555), .ZN(n580) );
  XOR2_X1 U434 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n367) );
  XNOR2_X1 U435 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n369) );
  XNOR2_X1 U438 ( .A(G134GAT), .B(G106GAT), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U440 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT79), .B(n401), .Z(n375) );
  NAND2_X1 U442 ( .A1(G232GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n382) );
  OR2_X1 U445 ( .A1(n580), .A2(n565), .ZN(n383) );
  OR2_X1 U446 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n391) );
  NOR2_X1 U448 ( .A1(n584), .A2(n555), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n387), .B(KEYINPUT45), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT68), .B(n546), .Z(n560) );
  INV_X1 U451 ( .A(n560), .ZN(n532) );
  NAND2_X1 U452 ( .A1(n388), .A2(n532), .ZN(n389) );
  NOR2_X1 U453 ( .A1(n577), .A2(n389), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n392), .B(KEYINPUT48), .ZN(n544) );
  XOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n394) );
  XNOR2_X1 U456 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U458 ( .A(KEYINPUT19), .B(n395), .ZN(n452) );
  XOR2_X1 U459 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n396) );
  XOR2_X1 U460 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U463 ( .A(n405), .B(n404), .Z(n407) );
  XNOR2_X1 U464 ( .A(G36GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n408) );
  NOR2_X1 U466 ( .A1(n544), .A2(n518), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT54), .ZN(n433) );
  XOR2_X1 U468 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n411) );
  XNOR2_X1 U469 ( .A(KEYINPUT1), .B(KEYINPUT95), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n424) );
  XOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT94), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT6), .B(KEYINPUT98), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U477 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U478 ( .A(G127GAT), .B(KEYINPUT0), .Z(n419) );
  XNOR2_X1 U479 ( .A(G113GAT), .B(G134GAT), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n447) );
  XNOR2_X1 U481 ( .A(n447), .B(n420), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n432) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(G120GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U488 ( .A(G29GAT), .B(G162GAT), .Z(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U491 ( .A(n432), .B(n431), .Z(n469) );
  INV_X1 U492 ( .A(n469), .ZN(n514) );
  NAND2_X1 U493 ( .A1(n433), .A2(n514), .ZN(n434) );
  INV_X1 U494 ( .A(n570), .ZN(n435) );
  NOR2_X1 U495 ( .A1(n470), .A2(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n454) );
  XOR2_X1 U498 ( .A(KEYINPUT86), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(G15GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT85), .B(G99GAT), .Z(n441) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(G190GAT), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U504 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(n446), .B(KEYINPUT65), .Z(n449) );
  XNOR2_X1 U508 ( .A(n447), .B(KEYINPUT20), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n453) );
  INV_X1 U511 ( .A(n455), .ZN(n549) );
  INV_X1 U512 ( .A(n549), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n566), .A2(n456), .ZN(n460) );
  XOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT123), .Z(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  NOR2_X1 U516 ( .A1(n577), .A2(n532), .ZN(n485) );
  NOR2_X1 U517 ( .A1(n528), .A2(n518), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT101), .B(n461), .Z(n462) );
  NOR2_X1 U519 ( .A1(n470), .A2(n462), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT25), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n528), .A2(n470), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT26), .B(n464), .Z(n569) );
  XOR2_X1 U523 ( .A(KEYINPUT27), .B(n518), .Z(n468) );
  NAND2_X1 U524 ( .A1(n569), .A2(n468), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n467), .A2(n514), .ZN(n473) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n543) );
  XOR2_X1 U528 ( .A(n470), .B(KEYINPUT28), .Z(n525) );
  INV_X1 U529 ( .A(n525), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n543), .A2(n471), .ZN(n530) );
  NAND2_X1 U531 ( .A1(n530), .A2(n528), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n473), .A2(n472), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n555), .A2(n482), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT107), .B(n474), .Z(n475) );
  NOR2_X1 U535 ( .A1(n584), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT37), .B(n476), .Z(n513) );
  NAND2_X1 U537 ( .A1(n485), .A2(n513), .ZN(n477) );
  NOR2_X1 U538 ( .A1(n500), .A2(n528), .ZN(n480) );
  INV_X1 U539 ( .A(G43GAT), .ZN(n478) );
  NOR2_X1 U540 ( .A1(n565), .A2(n555), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT16), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(n484), .Z(n503) );
  NAND2_X1 U544 ( .A1(n485), .A2(n503), .ZN(n495) );
  NOR2_X1 U545 ( .A1(n514), .A2(n495), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n518), .A2(n495), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(n489), .Z(n490) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n495), .A2(n528), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n492) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n525), .A2(n495), .ZN(n496) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n496), .Z(G1327GAT) );
  NOR2_X1 U559 ( .A1(n500), .A2(n514), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n500), .A2(n518), .ZN(n499) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U564 ( .A1(n525), .A2(n500), .ZN(n501) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NOR2_X1 U566 ( .A1(n549), .A2(n571), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(KEYINPUT108), .ZN(n512) );
  NAND2_X1 U568 ( .A1(n512), .A2(n503), .ZN(n508) );
  NOR2_X1 U569 ( .A1(n514), .A2(n508), .ZN(n504) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n518), .A2(n508), .ZN(n506) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n528), .A2(n508), .ZN(n507) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n525), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n514), .A2(n524), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n518), .A2(n524), .ZN(n519) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n528), .A2(n524), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT112), .B(n520), .Z(n521) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n523) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U594 ( .A(n527), .B(n526), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n544), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(n531), .ZN(n539) );
  NOR2_X1 U598 ( .A1(n539), .A2(n532), .ZN(n533) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n539), .A2(n549), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n539), .A2(n555), .ZN(n537) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n539), .A2(n558), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n545), .A2(n569), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n546), .A2(n557), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n557), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT52), .B(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n557), .ZN(n556) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n559), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n566), .A2(n580), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT124), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT125), .B(n564), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n583) );
  INV_X1 U637 ( .A(n583), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(n574), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U644 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

