//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  NAND2_X1  g000(.A1(G217), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT73), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n195), .C1(G119), .C2(new_n194), .ZN(new_n196));
  XNOR2_X1  g010(.A(G119), .B(G128), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT24), .B(G110), .Z(new_n198));
  OAI22_X1  g012(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(KEYINPUT74), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(G125), .A3(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n201), .B2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n198), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n205), .A2(new_n211), .A3(new_n207), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT75), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT75), .B1(new_n213), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT76), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(KEYINPUT77), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n217), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT75), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n226), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n217), .A3(new_n213), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n241), .B(new_n238), .C1(new_n227), .C2(new_n234), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n190), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n190), .A2(G902), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT78), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(new_n236), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n211), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G128), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n255), .A2(G137), .ZN(new_n258));
  OAI21_X1  g072(.A(G131), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n255), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .A4(new_n256), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n249), .B(new_n251), .C1(KEYINPUT1), .C2(new_n194), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n254), .A2(new_n259), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n263), .A3(new_n256), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(new_n265), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT0), .B(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n252), .A2(new_n278), .A3(KEYINPUT64), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n267), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G119), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT65), .B1(new_n192), .B2(G116), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n282), .A3(G119), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT2), .B(G113), .Z(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n269), .A2(new_n265), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(new_n274), .A3(new_n276), .A4(new_n279), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n287), .B(new_n288), .Z(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n267), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n248), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n281), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT28), .B1(new_n296), .B2(new_n293), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT26), .B(G101), .ZN(new_n299));
  INV_X1    g113(.A(G237), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n300), .A2(new_n221), .A3(G210), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n299), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n299), .A2(new_n301), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n301), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n298), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  INV_X1    g129(.A(new_n294), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n281), .A2(KEYINPUT30), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(new_n267), .C1(new_n270), .C2(new_n280), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n320), .B2(new_n289), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n315), .B1(new_n321), .B2(new_n309), .ZN(new_n322));
  INV_X1    g136(.A(new_n309), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n293), .B1(new_n317), .B2(new_n319), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT72), .B(new_n323), .C1(new_n324), .C2(new_n316), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n314), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n309), .A2(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g141(.A(G902), .B1(new_n298), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n313), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n295), .B2(new_n297), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n330), .B(KEYINPUT71), .C1(new_n295), .C2(new_n297), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n319), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n318), .B1(new_n292), .B2(new_n267), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n289), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n294), .A2(new_n309), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n338), .A2(new_n339), .A3(new_n343), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n294), .A2(new_n309), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n324), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT67), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT31), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(G472), .A2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(G472), .A2(new_n329), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n354), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n247), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G469), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n221), .A2(G227), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT80), .ZN(new_n362));
  XNOR2_X1  g176(.A(G110), .B(G140), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n366), .B2(G104), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G107), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n366), .A2(KEYINPUT3), .A3(G104), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n366), .B2(G104), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n367), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n369), .B2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(KEYINPUT3), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n367), .A4(new_n370), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n280), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n367), .A2(new_n370), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n383), .B2(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT82), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND4_X1   g200(.A1(KEYINPUT82), .A2(new_n373), .A3(new_n385), .A4(G101), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n381), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n254), .A2(new_n266), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n369), .A2(G107), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n366), .A2(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(G101), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n380), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n380), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT10), .B(new_n390), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n380), .A2(new_n394), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n291), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n388), .A2(new_n397), .A3(new_n270), .A4(new_n400), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n365), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND4_X1   g218(.A1(new_n380), .A2(new_n394), .A3(new_n266), .A4(new_n254), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n380), .A2(new_n394), .B1(new_n254), .B2(new_n266), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n291), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT12), .B(new_n291), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(new_n403), .A3(new_n365), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n360), .B(new_n237), .C1(new_n404), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(G469), .A2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n403), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n364), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n403), .A3(new_n365), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(G469), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n420), .B2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT79), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(KEYINPUT84), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n283), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G113), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n430), .A2(new_n434), .B1(new_n287), .B2(new_n288), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n395), .B2(new_n396), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n386), .A2(new_n387), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n381), .A2(new_n289), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n436), .B(new_n440), .C1(new_n437), .C2(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n439), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n280), .A2(G125), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n389), .A2(new_n201), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G224), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n440), .B(KEYINPUT8), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n380), .A2(KEYINPUT86), .A3(new_n394), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n380), .A2(new_n457), .A3(new_n394), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n460), .B2(new_n435), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n287), .A2(new_n288), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n431), .B(new_n283), .C1(new_n286), .C2(new_n284), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n433), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n459), .B2(new_n458), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n455), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n451), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n447), .A2(new_n448), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n447), .B2(new_n448), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n471), .A3(new_n443), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n472), .A2(new_n237), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n453), .A2(new_n454), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n454), .B1(new_n453), .B2(new_n473), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n429), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G237), .A2(G953), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n477), .A2(G143), .A3(G214), .ZN(new_n478));
  AOI21_X1  g292(.A(G143), .B1(new_n477), .B2(G214), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n300), .A2(new_n221), .A3(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n250), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(G143), .A3(G214), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n264), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT19), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n210), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n202), .A2(KEYINPUT19), .A3(new_n204), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n211), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n485), .A2(new_n209), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n482), .A2(new_n483), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(KEYINPUT87), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  INV_X1    g308(.A(new_n491), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n482), .A2(new_n494), .A3(new_n495), .A4(new_n483), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n202), .A2(G146), .A3(new_n204), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n493), .A2(new_n496), .B1(new_n212), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT88), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n212), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n485), .A2(new_n209), .A3(new_n489), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n369), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT89), .B1(new_n480), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n492), .A2(new_n512), .A3(KEYINPUT17), .A4(G131), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n480), .A2(new_n510), .A3(new_n484), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n215), .A2(new_n216), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n480), .A2(new_n484), .A3(KEYINPUT90), .A4(new_n510), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n507), .A3(new_n502), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT20), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n507), .A3(new_n502), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n507), .B1(new_n520), .B2(new_n502), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n237), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT91), .B(new_n237), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(G475), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(G234), .A2(G237), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n536), .A2(G952), .A3(new_n221), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT21), .B(G898), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(G902), .A3(G953), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n282), .A2(G122), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n282), .B2(G122), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n282), .A3(G122), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n543), .A2(new_n545), .B1(new_n546), .B2(KEYINPUT92), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n366), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G122), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G116), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n551), .A3(new_n366), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n250), .A2(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n194), .A2(G143), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n255), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n255), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n552), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n366), .B1(new_n543), .B2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n194), .B2(G143), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n250), .A2(KEYINPUT13), .A3(G128), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(G134), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n549), .A2(new_n558), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n420), .A2(new_n188), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI221_X1 g384(.A(new_n568), .B1(new_n561), .B2(new_n566), .C1(new_n549), .C2(new_n558), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT93), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n567), .A2(new_n573), .A3(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n237), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G478), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(KEYINPUT15), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n575), .B(new_n577), .Z(new_n578));
  NAND4_X1  g392(.A1(new_n528), .A2(new_n535), .A3(new_n542), .A4(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n476), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n359), .A2(new_n428), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n351), .B2(new_n237), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n348), .A2(new_n349), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n585), .A2(KEYINPUT31), .B1(new_n333), .B2(new_n334), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n353), .B1(new_n586), .B2(new_n345), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n247), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n429), .B(new_n542), .C1(new_n474), .C2(new_n475), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n534), .A2(G475), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n592), .A2(new_n533), .B1(new_n525), .B2(new_n527), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT33), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n572), .A2(new_n596), .A3(new_n574), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n572), .A2(new_n599), .A3(new_n596), .A4(new_n574), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n595), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n576), .A2(G902), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(new_n576), .B2(new_n575), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n591), .B1(new_n593), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n528), .A2(new_n535), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n598), .A2(new_n600), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n594), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n575), .A2(new_n576), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n605), .A2(KEYINPUT95), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  AND4_X1   g425(.A1(new_n428), .A2(new_n588), .A3(new_n590), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(new_n578), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n589), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n588), .A2(new_n428), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  AOI21_X1  g434(.A(KEYINPUT77), .B1(new_n220), .B2(new_n226), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n218), .A2(new_n219), .A3(new_n233), .A4(new_n225), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n239), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n241), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n239), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n220), .B(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n626), .A2(new_n190), .B1(new_n245), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(new_n584), .A3(new_n587), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n428), .A3(new_n580), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  NAND2_X1  g447(.A1(new_n356), .A2(new_n358), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n629), .A2(new_n476), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n616), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n541), .A2(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n538), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n403), .A2(new_n365), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n640), .A2(new_n402), .B1(new_n415), .B2(new_n364), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n641), .B2(G902), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n425), .B(new_n422), .C1(new_n642), .C2(new_n413), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT84), .B1(new_n419), .B2(new_n423), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n637), .B(new_n639), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT96), .B1(new_n636), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n593), .A2(new_n615), .A3(new_n639), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n426), .B2(new_n427), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n634), .A4(new_n635), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XNOR2_X1  g466(.A(new_n639), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n428), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n290), .A2(new_n294), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n585), .B1(new_n657), .B2(new_n313), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n583), .B1(new_n658), .B2(new_n237), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n351), .B2(new_n355), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n660), .A2(new_n358), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n474), .A2(new_n475), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT38), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n578), .B1(new_n528), .B2(new_n535), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n629), .A2(new_n429), .A3(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n655), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(new_n636), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n605), .A2(new_n609), .A3(new_n639), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n426), .B2(new_n427), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT97), .B(G146), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G48));
  OAI21_X1  g489(.A(new_n237), .B1(new_n404), .B2(new_n412), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n421), .A3(new_n413), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n359), .A2(new_n590), .A3(new_n611), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT98), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G15));
  NAND3_X1  g497(.A1(new_n359), .A2(new_n617), .A3(new_n679), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NOR2_X1   g499(.A1(new_n678), .A2(new_n579), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n634), .A2(new_n635), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NAND2_X1  g502(.A1(new_n351), .A2(new_n237), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n350), .A2(KEYINPUT99), .A3(new_n331), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n345), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT99), .B1(new_n350), .B2(new_n331), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n352), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n605), .A2(new_n615), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n589), .A2(new_n696), .A3(new_n678), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n243), .A2(new_n246), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NOR2_X1   g514(.A1(new_n476), .A2(new_n678), .ZN(new_n701));
  INV_X1    g515(.A(new_n671), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n628), .A2(new_n245), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n243), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n690), .A2(new_n705), .A3(new_n694), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n201), .ZN(G27));
  NAND2_X1  g522(.A1(new_n329), .A2(G472), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n351), .A2(new_n355), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT32), .B1(new_n351), .B2(new_n352), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n698), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT100), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n634), .A2(new_n715), .A3(new_n698), .ZN(new_n716));
  INV_X1    g530(.A(new_n429), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n474), .A2(new_n475), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n421), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n642), .B2(new_n413), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n528), .A2(new_n535), .B1(new_n607), .B2(new_n608), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n639), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n716), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n419), .A2(new_n421), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n453), .A2(new_n473), .ZN(new_n727));
  INV_X1    g541(.A(new_n454), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n453), .A2(new_n454), .A3(new_n473), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n429), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n634), .A2(new_n732), .A3(new_n702), .A4(new_n698), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n723), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n725), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n725), .A2(KEYINPUT101), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n264), .ZN(G33));
  NAND4_X1  g554(.A1(new_n359), .A2(new_n637), .A3(new_n639), .A4(new_n732), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  XNOR2_X1  g556(.A(new_n718), .B(KEYINPUT103), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n593), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n605), .A2(KEYINPUT102), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT43), .A4(new_n609), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n605), .B2(new_n603), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(new_n705), .C1(new_n587), .C2(new_n584), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n743), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n751), .A2(new_n752), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n641), .A2(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n416), .A2(new_n417), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n761), .A3(G469), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n414), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n413), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n421), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n653), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT105), .B(G137), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT47), .B(new_n421), .C1(new_n766), .C2(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n634), .A2(new_n698), .A3(new_n731), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n702), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  AND2_X1   g594(.A1(new_n695), .A2(new_n698), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n538), .B1(new_n747), .B2(new_n749), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n678), .A2(KEYINPUT111), .A3(new_n429), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT111), .B1(new_n678), .B2(new_n429), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n663), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n781), .A2(new_n782), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n785), .B1(new_n792), .B2(new_n789), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n677), .A2(new_n413), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n423), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n743), .B(new_n783), .C1(new_n777), .C2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n690), .A2(new_n705), .A3(new_n694), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n731), .A2(new_n678), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n782), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n731), .A2(new_n678), .A3(new_n538), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n605), .A2(new_n609), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n661), .A2(new_n803), .A3(new_n698), .A4(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n794), .A2(new_n799), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n661), .A2(new_n803), .A3(new_n698), .A4(new_n611), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(G952), .A3(new_n221), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n714), .A2(new_n716), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n782), .A4(new_n801), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n782), .A2(new_n801), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT48), .B1(new_n813), .B2(new_n809), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n808), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n781), .A2(new_n701), .A3(new_n782), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n815), .A2(KEYINPUT116), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n815), .B2(new_n818), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n806), .A2(KEYINPUT51), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n802), .A2(new_n805), .A3(KEYINPUT113), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n802), .B2(new_n805), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n794), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n794), .B(KEYINPUT114), .C1(new_n824), .C2(new_n823), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n611), .A2(new_n590), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n698), .B(new_n679), .C1(new_n711), .C2(new_n712), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n580), .B1(new_n644), .B2(new_n643), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n584), .A2(new_n587), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n705), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n687), .B1(new_n833), .B2(new_n713), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n616), .B1(new_n593), .B2(new_n603), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n588), .A2(new_n428), .A3(new_n590), .A4(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n840), .A2(new_n699), .A3(new_n684), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n671), .A2(new_n726), .A3(new_n731), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n800), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT106), .B1(new_n706), .B2(new_n722), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n629), .A2(new_n731), .ZN(new_n847));
  INV_X1    g661(.A(new_n639), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n605), .A2(new_n615), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n428), .A2(new_n847), .A3(new_n634), .A4(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n741), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n838), .A2(new_n841), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT107), .B1(new_n739), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n725), .A2(KEYINPUT101), .A3(new_n734), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT101), .B1(new_n725), .B2(new_n734), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n842), .B1(new_n800), .B2(new_n843), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n706), .A2(new_n722), .A3(KEYINPUT106), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n741), .B(new_n850), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(new_n699), .A3(new_n684), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n680), .A2(new_n581), .A3(new_n631), .A4(new_n687), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT107), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n707), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n664), .B(new_n429), .C1(new_n475), .C2(new_n474), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n660), .B2(new_n358), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n705), .A2(new_n726), .A3(new_n848), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n670), .A2(new_n672), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n651), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n651), .A2(new_n869), .A3(KEYINPUT52), .A4(new_n865), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n853), .A2(new_n864), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(KEYINPUT109), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n869), .A2(KEYINPUT52), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT108), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n651), .B2(new_n865), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT108), .B(new_n707), .C1(new_n646), .C2(new_n650), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT109), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n870), .A2(new_n884), .A3(new_n871), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n877), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n862), .A2(KEYINPUT53), .A3(new_n735), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n875), .A2(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(new_n876), .A3(new_n864), .A4(new_n853), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n830), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(G952), .A2(G953), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n663), .A2(new_n746), .A3(new_n745), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n609), .A2(new_n423), .A3(new_n429), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n698), .A3(new_n661), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n896), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n221), .A2(G952), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT120), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n888), .A2(new_n237), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n444), .A2(new_n446), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n452), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n909), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n875), .A2(new_n876), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n886), .A2(new_n887), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n921), .A3(G902), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT118), .B1(new_n888), .B2(new_n237), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n728), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n923), .A3(new_n728), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT119), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n915), .B1(new_n926), .B2(new_n928), .ZN(G51));
  NAND2_X1  g743(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n931), .A3(new_n890), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n920), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n414), .B(KEYINPUT57), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n404), .A2(new_n412), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n762), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n922), .A2(new_n923), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n908), .B1(new_n937), .B2(new_n939), .ZN(G54));
  AND2_X1   g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n922), .A2(new_n923), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n522), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n942), .A2(KEYINPUT122), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT122), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n922), .A2(new_n923), .A3(new_n522), .A4(new_n941), .ZN(new_n946));
  INV_X1    g760(.A(new_n908), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(G60));
  XNOR2_X1  g763(.A(new_n601), .B(KEYINPUT123), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT59), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n933), .A2(new_n932), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n890), .B2(new_n893), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n909), .B1(new_n955), .B2(new_n950), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G63));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n187), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n888), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(new_n628), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n235), .A2(new_n236), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT125), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n909), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n959), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n958), .A2(new_n920), .A3(new_n628), .A4(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n960), .A2(new_n963), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n960), .A2(new_n628), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n972), .B(new_n973), .C1(new_n968), .C2(new_n969), .ZN(new_n974));
  OAI22_X1  g788(.A1(new_n967), .A2(KEYINPUT61), .B1(new_n971), .B2(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n539), .B2(new_n450), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n861), .A2(new_n860), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n912), .B1(G898), .B2(new_n221), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  NAND2_X1  g794(.A1(new_n487), .A2(new_n488), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n320), .B(new_n981), .Z(new_n982));
  OR2_X1    g796(.A1(new_n881), .A2(new_n882), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n668), .A3(new_n673), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g800(.A(new_n654), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(new_n359), .A3(new_n718), .A4(new_n839), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n771), .A2(new_n779), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n982), .B1(new_n990), .B2(new_n221), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n809), .A2(new_n866), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n770), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n856), .A2(new_n741), .A3(new_n779), .A4(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n994), .A2(new_n673), .A3(new_n771), .A4(new_n983), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(G953), .ZN(new_n996));
  INV_X1    g810(.A(G900), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n982), .B1(new_n997), .B2(new_n221), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(G227), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n1001), .B2(new_n997), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  INV_X1    g819(.A(new_n977), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n990), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n321), .A2(new_n323), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1007), .A2(KEYINPUT127), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(KEYINPUT127), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n995), .B2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n323), .A3(new_n321), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n585), .A2(new_n322), .A3(new_n325), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n891), .A2(new_n892), .A3(new_n1005), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1012), .A2(new_n947), .A3(new_n1014), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1009), .A2(new_n1010), .A3(new_n1015), .ZN(G57));
endmodule


