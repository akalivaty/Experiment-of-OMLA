//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT72), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(G64gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT71), .ZN(new_n214));
  NAND2_X1  g013(.A1(G226gat), .A2(G233gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(KEYINPUT66), .B2(KEYINPUT24), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n227), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT23), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n219), .B(KEYINPUT65), .C1(new_n220), .C2(new_n221), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n224), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n236));
  AND2_X1   g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n226), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT28), .ZN(new_n245));
  OR3_X1    g044(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(new_n226), .C1(new_n237), .C2(new_n238), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n251), .A3(new_n229), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  INV_X1    g054(.A(new_n229), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT24), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n228), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(new_n233), .A3(new_n224), .A4(new_n234), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n254), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n216), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n241), .A2(KEYINPUT67), .A3(new_n242), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n250), .B1(new_n267), .B2(new_n226), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n222), .A2(new_n223), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n233), .A3(new_n234), .A4(new_n247), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n268), .A2(new_n252), .B1(new_n270), .B2(new_n259), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n215), .B1(new_n272), .B2(new_n236), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n214), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT29), .B1(new_n272), .B2(new_n236), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n275), .B2(new_n216), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n213), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n216), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n213), .B(new_n278), .C1(new_n275), .C2(new_n216), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT30), .B(new_n205), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n263), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n214), .B1(new_n284), .B2(new_n215), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n275), .B2(new_n216), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(new_n214), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n279), .B1(new_n287), .B2(new_n213), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n205), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n277), .A2(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(new_n205), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G141gat), .B(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(KEYINPUT2), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n305), .B(KEYINPUT74), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT1), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT68), .B(G120gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n313), .B(new_n315), .C1(new_n318), .C2(new_n311), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT76), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G162gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n325), .A3(G155gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n327));
  INV_X1    g126(.A(new_n305), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n328), .A2(new_n307), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n330));
  INV_X1    g129(.A(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT75), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n327), .B(new_n329), .C1(new_n330), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n333), .A2(G148gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n331), .A2(G141gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT75), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n342), .A2(new_n343), .B1(new_n326), .B2(KEYINPUT2), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT77), .B1(new_n344), .B2(new_n329), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n310), .B(new_n321), .C1(new_n338), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n336), .A2(new_n337), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT77), .A3(new_n329), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n309), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n321), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n310), .B1(new_n338), .B2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT3), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n320), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n350), .B2(new_n321), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n320), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n359), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n354), .A2(KEYINPUT78), .A3(new_n320), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n360), .A2(new_n366), .A3(KEYINPUT5), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n360), .A2(new_n366), .A3(new_n369), .A4(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n352), .A2(KEYINPUT81), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n350), .A2(new_n373), .A3(new_n351), .A4(new_n321), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n347), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n364), .A2(KEYINPUT5), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n375), .A2(new_n358), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n303), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n302), .B(new_n377), .C1(new_n368), .C2(new_n370), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT6), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n378), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n302), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n297), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT82), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n321), .B1(new_n387), .B2(new_n271), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n236), .A2(new_n254), .A3(new_n320), .A4(new_n261), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G227gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT34), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n388), .B2(new_n389), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT69), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n388), .A2(new_n393), .A3(new_n389), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G71gat), .ZN(new_n405));
  INV_X1    g204(.A(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n402), .B(KEYINPUT32), .C1(new_n403), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(KEYINPUT32), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n402), .A2(new_n403), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n398), .A2(new_n399), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n401), .A2(new_n409), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n409), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n413), .A3(new_n400), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OR3_X1    g218(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n212), .B1(new_n357), .B2(new_n263), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n212), .B2(new_n263), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n350), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G228gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n392), .ZN(new_n430));
  AOI211_X1 g229(.A(KEYINPUT3), .B(new_n309), .C1(new_n348), .C2(new_n349), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n213), .B1(new_n431), .B2(KEYINPUT29), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT85), .B1(new_n350), .B2(new_n426), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n428), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT84), .B1(new_n425), .B2(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(new_n430), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G22gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(new_n440), .A3(G22gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445));
  INV_X1    g244(.A(G50gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n443), .B(new_n444), .C1(KEYINPUT86), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n444), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  AOI21_X1  g252(.A(G22gat), .B1(new_n437), .B2(new_n440), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n452), .B(new_n449), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n414), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n416), .A2(new_n417), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT36), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n423), .A2(new_n451), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n449), .B1(new_n454), .B2(new_n453), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n443), .B2(new_n444), .ZN(new_n462));
  INV_X1    g261(.A(new_n451), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT35), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n382), .A2(new_n302), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n377), .B1(new_n368), .B2(new_n370), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT6), .B1(new_n467), .B2(new_n303), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n383), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n297), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n386), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n451), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n419), .A2(KEYINPUT89), .A3(new_n420), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT89), .B1(new_n419), .B2(new_n420), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(new_n385), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n363), .A2(new_n365), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n359), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n375), .A2(new_n358), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT39), .B(new_n481), .C1(new_n482), .C2(new_n359), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n359), .B1(new_n375), .B2(new_n358), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT39), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n302), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n483), .A2(KEYINPUT40), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT40), .B1(new_n483), .B2(new_n486), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n296), .A2(new_n489), .A3(new_n466), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n274), .A2(new_n213), .A3(new_n276), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n286), .A2(new_n212), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT37), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n491), .A2(new_n495), .A3(KEYINPUT37), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n288), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n499), .C1(new_n277), .C2(new_n280), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n497), .B(new_n293), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT38), .B1(new_n288), .B2(new_n205), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n279), .B(KEYINPUT37), .C1(new_n287), .C2(new_n213), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT38), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT88), .B1(new_n292), .B2(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n503), .A2(new_n504), .B1(new_n508), .B2(new_n293), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n490), .B1(new_n470), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n423), .A2(new_n458), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n475), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n473), .A2(new_n479), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G197gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT11), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n217), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G15gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n442), .ZN(new_n521));
  NAND2_X1  g320(.A1(G15gat), .A2(G22gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n526), .A3(new_n522), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT93), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(G8gat), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n523), .B(KEYINPUT94), .C1(new_n524), .C2(G1gat), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n527), .A4(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G43gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(G50gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n446), .A2(G43gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT90), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  INV_X1    g340(.A(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n446), .A2(G43gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n537), .A2(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n540), .A2(new_n547), .A3(KEYINPUT15), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n538), .B2(new_n539), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n543), .A2(new_n545), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n543), .B2(new_n545), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n546), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n551), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n552), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT92), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n552), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n536), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n565), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n568), .B2(new_n536), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT18), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n519), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n571), .B(new_n564), .C1(new_n568), .C2(new_n536), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n530), .A2(new_n535), .ZN(new_n577));
  INV_X1    g376(.A(new_n563), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n543), .A2(new_n545), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT91), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n543), .A2(new_n545), .A3(new_n555), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n551), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n546), .A4(new_n554), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n562), .B1(new_n584), .B2(new_n552), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n536), .A2(new_n561), .A3(new_n563), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n571), .B(KEYINPUT13), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n590), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT18), .A2(new_n576), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n536), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n572), .A3(new_n586), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT18), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n576), .A2(KEYINPUT18), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n594), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n519), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n513), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G183gat), .B(G211gat), .Z(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT99), .B(KEYINPUT20), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(G57gat), .A2(G64gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G57gat), .A2(G64gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G71gat), .B(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n536), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT101), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n631), .A2(new_n632), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n627), .A3(new_n633), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n636), .B2(new_n640), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n613), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n634), .A2(new_n635), .A3(new_n628), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n627), .B1(new_n639), .B2(new_n633), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n637), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n641), .A3(new_n612), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT7), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT7), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n652), .A2(KEYINPUT103), .A3(G85gat), .A4(G92gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G99gat), .B(G106gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  INV_X1    g455(.A(G85gat), .ZN(new_n657));
  INV_X1    g456(.A(G92gat), .ZN(new_n658));
  AOI22_X1  g457(.A1(KEYINPUT8), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n654), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n654), .B2(new_n659), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n568), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n578), .B2(new_n585), .ZN(new_n664));
  NAND3_X1  g463(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667));
  XOR2_X1   g466(.A(G190gat), .B(G218gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n667), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT102), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G134gat), .B(G162gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n670), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n649), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n607), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n654), .A2(new_n659), .ZN(new_n681));
  INV_X1    g480(.A(new_n655), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n654), .A2(new_n655), .A3(new_n659), .ZN(new_n684));
  INV_X1    g483(.A(new_n625), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n624), .B(new_n625), .C1(new_n660), .C2(new_n661), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n663), .A2(new_n626), .A3(KEYINPUT10), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n680), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n680), .B1(new_n687), .B2(new_n688), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(G120gat), .B(G148gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n218), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(G204gat), .Z(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n695), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n680), .B(KEYINPUT107), .Z(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n690), .B2(new_n692), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n700), .B1(new_n706), .B2(new_n696), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n702), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n679), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n470), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n526), .ZN(G1324gat));
  NOR2_X1   g513(.A1(new_n524), .A2(new_n533), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n712), .A2(new_n297), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n524), .A2(new_n533), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n712), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n296), .ZN(new_n722));
  AOI22_X1  g521(.A1(G8gat), .A2(new_n722), .B1(new_n716), .B2(new_n717), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n723), .B2(new_n719), .ZN(G1325gat));
  NOR3_X1   g523(.A1(new_n712), .A2(new_n520), .A3(new_n511), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n476), .A2(new_n477), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n520), .B2(new_n728), .ZN(G1326gat));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n475), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT43), .B(G22gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1327gat));
  INV_X1    g531(.A(new_n649), .ZN(new_n733));
  INV_X1    g532(.A(new_n677), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n733), .A2(new_n710), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n607), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n470), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n541), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n733), .A2(new_n710), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n513), .A2(new_n743), .A3(new_n677), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n513), .B2(new_n677), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n606), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n470), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n741), .A2(new_n747), .ZN(G1328gat));
  NAND3_X1  g547(.A1(new_n738), .A2(new_n542), .A3(new_n296), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT46), .Z(new_n750));
  OAI21_X1  g549(.A(G36gat), .B1(new_n746), .B2(new_n297), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n607), .A2(new_n537), .A3(new_n736), .A4(new_n737), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n726), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT110), .B1(new_n753), .B2(new_n726), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G43gat), .B1(new_n746), .B2(new_n511), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1330gat));
  OAI21_X1  g561(.A(G50gat), .B1(new_n746), .B2(new_n475), .ZN(new_n763));
  INV_X1    g562(.A(new_n475), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n738), .A2(new_n446), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g566(.A(new_n678), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n606), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n513), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n710), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n739), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n296), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  INV_X1    g578(.A(new_n511), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G71gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  INV_X1    g582(.A(G71gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n726), .A2(new_n711), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n783), .B1(new_n782), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT50), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n771), .A2(new_n764), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n470), .A2(G85gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n733), .A2(new_n606), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n513), .A2(new_n677), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT113), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n710), .B(new_n797), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n710), .B(new_n799), .C1(new_n744), .C2(new_n745), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT112), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n739), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n809), .B2(new_n657), .ZN(G1336gat));
  NOR3_X1   g609(.A1(new_n297), .A2(G92gat), .A3(new_n711), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n804), .B2(new_n805), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(G92gat), .B1(new_n807), .B2(new_n297), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n811), .B(KEYINPUT114), .Z(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n802), .B2(new_n803), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  INV_X1    g617(.A(new_n799), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n513), .A2(new_n677), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT44), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n513), .A2(new_n743), .A3(new_n677), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n823), .B2(new_n710), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n296), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n817), .B1(new_n826), .B2(G92gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n815), .B1(new_n827), .B2(new_n813), .ZN(G1337gat));
  AND2_X1   g627(.A1(new_n808), .A2(new_n780), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n804), .A2(new_n805), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n785), .A2(new_n406), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n829), .A2(new_n406), .B1(new_n830), .B2(new_n831), .ZN(G1338gat));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(G106gat), .B1(new_n807), .B2(new_n475), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n475), .A2(G106gat), .A3(new_n711), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n833), .B(new_n834), .C1(new_n830), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n802), .B2(new_n803), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n764), .B1(new_n824), .B2(new_n825), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(G106gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n840), .B2(new_n833), .ZN(G1339gat));
  AOI21_X1  g640(.A(KEYINPUT96), .B1(new_n588), .B2(new_n590), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n592), .B(new_n589), .C1(new_n586), .C2(new_n587), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n597), .A2(new_n598), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n574), .B1(new_n597), .B2(new_n598), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n846), .A2(new_n575), .B1(new_n604), .B2(new_n519), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n678), .A2(new_n711), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n702), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n701), .B1(new_n706), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n680), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n690), .A2(new_n692), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT106), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n690), .A2(new_n692), .A3(new_n691), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n690), .A2(new_n692), .A3(new_n705), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  INV_X1    g659(.A(new_n858), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n695), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n851), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT55), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(new_n856), .B2(new_n858), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n695), .A2(new_n860), .A3(new_n861), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n851), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n849), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n517), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n569), .A2(new_n572), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n846), .B2(new_n575), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n677), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n870), .A2(new_n606), .B1(new_n875), .B2(new_n710), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT116), .B(new_n876), .C1(new_n877), .C2(new_n677), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n649), .ZN(new_n879));
  INV_X1    g678(.A(new_n874), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n601), .A2(new_n710), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n867), .A2(new_n868), .A3(new_n851), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n868), .B1(new_n867), .B2(new_n851), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n702), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(new_n847), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n734), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT116), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n848), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n848), .B(KEYINPUT117), .C1(new_n879), .C2(new_n887), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n475), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n470), .A2(new_n296), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n890), .A2(new_n895), .A3(new_n475), .A4(new_n891), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n893), .A2(new_n727), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G113gat), .B1(new_n897), .B2(new_n847), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n890), .A2(new_n891), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n475), .A2(new_n460), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n739), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n901), .A2(KEYINPUT120), .A3(new_n739), .A4(new_n902), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n296), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n311), .A3(new_n606), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n900), .A2(new_n908), .ZN(G1340gat));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n318), .A3(new_n710), .ZN(new_n910));
  OAI21_X1  g709(.A(G120gat), .B1(new_n897), .B2(new_n711), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1341gat));
  INV_X1    g711(.A(G127gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n913), .A3(new_n649), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n907), .A2(new_n733), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n913), .ZN(G1342gat));
  INV_X1    g715(.A(G134gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n907), .A2(new_n917), .A3(new_n677), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n919));
  OAI21_X1  g718(.A(G134gat), .B1(new_n897), .B2(new_n734), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n907), .A2(new_n921), .A3(new_n917), .A4(new_n677), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G1343gat));
  INV_X1    g722(.A(KEYINPUT57), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n901), .A2(new_n924), .A3(new_n764), .ZN(new_n925));
  INV_X1    g724(.A(new_n848), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n886), .B(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n876), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n649), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT57), .B1(new_n929), .B2(new_n475), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n894), .A2(new_n511), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n925), .A2(new_n930), .A3(new_n606), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G141gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n901), .A2(new_n739), .ZN(new_n935));
  INV_X1    g734(.A(new_n459), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n847), .A2(G141gat), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n935), .A2(new_n297), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n939), .A3(KEYINPUT58), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT58), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n933), .B(new_n938), .C1(KEYINPUT122), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1344gat));
  NAND3_X1  g742(.A1(new_n935), .A2(new_n297), .A3(new_n936), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n331), .A3(new_n710), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n925), .A2(new_n931), .A3(new_n930), .ZN(new_n947));
  AOI211_X1 g746(.A(KEYINPUT59), .B(new_n331), .C1(new_n947), .C2(new_n710), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n901), .A2(new_n764), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT57), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n733), .B1(new_n886), .B2(new_n876), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n924), .B(new_n764), .C1(new_n926), .C2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n951), .A2(new_n710), .A3(new_n931), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n954), .B2(G148gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n946), .B1(new_n948), .B2(new_n955), .ZN(G1345gat));
  INV_X1    g755(.A(G155gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n944), .B2(new_n649), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n649), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1346gat));
  NAND2_X1  g764(.A1(new_n947), .A2(new_n677), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n323), .A2(new_n325), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n947), .A2(KEYINPUT124), .A3(new_n677), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n945), .A2(new_n969), .A3(new_n677), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1347gat));
  NOR2_X1   g773(.A1(new_n739), .A2(new_n297), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n893), .A2(new_n727), .A3(new_n896), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G169gat), .B1(new_n976), .B2(new_n847), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n901), .A2(new_n902), .A3(new_n975), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(new_n217), .A3(new_n606), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT125), .ZN(G1348gat));
  NOR3_X1   g780(.A1(new_n976), .A2(new_n218), .A3(new_n711), .ZN(new_n982));
  AOI21_X1  g781(.A(G176gat), .B1(new_n978), .B2(new_n710), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(G1349gat));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n985), .A2(KEYINPUT60), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n985), .A2(KEYINPUT60), .ZN(new_n987));
  OAI21_X1  g786(.A(G183gat), .B1(new_n976), .B2(new_n649), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n978), .A2(new_n267), .A3(new_n733), .ZN(new_n989));
  AOI211_X1 g788(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  AND4_X1   g789(.A1(new_n985), .A2(new_n988), .A3(KEYINPUT60), .A4(new_n989), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(G1350gat));
  OAI21_X1  g791(.A(G190gat), .B1(new_n976), .B2(new_n734), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT61), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n226), .A3(new_n677), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1351gat));
  AND2_X1   g795(.A1(new_n951), .A2(new_n953), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n780), .A2(new_n739), .A3(new_n297), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n606), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G197gat), .ZN(new_n1000));
  INV_X1    g799(.A(new_n950), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(new_n998), .ZN(new_n1002));
  OR2_X1    g801(.A1(new_n847), .A2(G197gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1352gat));
  NAND3_X1  g803(.A1(new_n997), .A2(new_n710), .A3(new_n998), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(G204gat), .ZN(new_n1006));
  OR4_X1    g805(.A1(KEYINPUT62), .A2(new_n1002), .A3(G204gat), .A4(new_n711), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n1001), .A2(new_n998), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(new_n710), .ZN(new_n1009));
  OAI21_X1  g808(.A(KEYINPUT62), .B1(new_n1009), .B2(G204gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(G1353gat));
  NAND3_X1  g810(.A1(new_n1008), .A2(new_n207), .A3(new_n733), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n951), .A2(new_n733), .A3(new_n953), .A4(new_n998), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  OAI21_X1  g815(.A(new_n208), .B1(new_n1002), .B2(new_n734), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n734), .A2(new_n208), .ZN(new_n1018));
  NAND4_X1  g817(.A1(new_n951), .A2(new_n953), .A3(new_n998), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1017), .A2(new_n1022), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1021), .A2(new_n1023), .ZN(G1355gat));
endmodule


