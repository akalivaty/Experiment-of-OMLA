//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(new_n194), .C1(G119), .C2(new_n193), .ZN(new_n195));
  XNOR2_X1  g009(.A(G119), .B(G128), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT24), .B(G110), .Z(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT16), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n206), .A3(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(new_n202), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n198), .B(new_n207), .C1(G146), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n206), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n207), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n217), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n209), .A2(new_n215), .A3(new_n220), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n224), .B2(new_n188), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n189), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n189), .A2(G902), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n191), .B2(G116), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n233), .A3(G119), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n211), .A2(G143), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n243), .A2(KEYINPUT65), .A3(G146), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT65), .B1(new_n243), .B2(G146), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n241), .B(new_n242), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT11), .A3(G134), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(G137), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n254), .A2(G137), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n256), .A2(G134), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n261), .B(G131), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G134), .B(G137), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT66), .B1(new_n265), .B2(new_n258), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n252), .A2(new_n260), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n259), .A3(new_n257), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n260), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n243), .A2(G146), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n211), .B2(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n243), .A2(KEYINPUT65), .A3(G146), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n241), .B2(new_n249), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT0), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n193), .A3(KEYINPUT64), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(KEYINPUT0), .B2(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n276), .A2(new_n277), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n267), .A2(new_n268), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n268), .B1(new_n267), .B2(new_n285), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT68), .B(new_n240), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n240), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n271), .A2(new_n284), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n266), .A2(new_n260), .A3(new_n264), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n276), .A2(new_n242), .B1(new_n248), .B2(new_n250), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT30), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n267), .A2(new_n268), .A3(new_n285), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n267), .A3(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n288), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n302));
  NOR2_X1   g116(.A1(G237), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G210), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n302), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G101), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n300), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n297), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n240), .B1(new_n290), .B2(new_n293), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n313), .B2(new_n297), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n307), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n240), .B1(new_n286), .B2(new_n287), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n290), .A2(new_n293), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT68), .B1(new_n320), .B2(new_n289), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n318), .B(new_n307), .C1(new_n322), .C2(new_n288), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT70), .B1(new_n300), .B2(new_n308), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n317), .B1(new_n325), .B2(KEYINPUT31), .ZN(new_n326));
  NOR2_X1   g140(.A1(G472), .A2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT32), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n294), .A2(new_n295), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n299), .B1(new_n330), .B2(new_n240), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n298), .B(new_n289), .C1(new_n294), .C2(new_n295), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n308), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n318), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n309), .A2(new_n316), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n327), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n311), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(KEYINPUT29), .A3(new_n308), .A4(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n300), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n307), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n315), .B2(new_n307), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n348), .B(new_n188), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G472), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n232), .B1(new_n341), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G469), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n188), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT73), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(G104), .ZN(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n367), .B2(new_n369), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n375), .A2(new_n376), .A3(new_n252), .ZN(new_n377));
  INV_X1    g191(.A(new_n246), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n193), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n276), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n372), .A2(new_n374), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n271), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT12), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(KEYINPUT12), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n252), .A2(KEYINPUT10), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n375), .B2(new_n376), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n381), .B2(new_n382), .ZN(new_n393));
  INV_X1    g207(.A(new_n271), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n369), .B1(new_n360), .B2(new_n362), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n368), .A2(G107), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n396), .A2(new_n365), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n372), .A3(KEYINPUT4), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(G101), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n284), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n391), .A2(new_n393), .A3(new_n394), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G140), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n218), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n271), .B(new_n386), .C1(new_n377), .C2(new_n383), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n389), .A2(new_n403), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n391), .A2(new_n393), .A3(new_n402), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n271), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n403), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n406), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n358), .B1(new_n414), .B2(new_n357), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n382), .A2(KEYINPUT75), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n292), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n381), .A2(new_n382), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n394), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n387), .A2(new_n388), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n408), .B(new_n403), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n406), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n411), .A2(new_n403), .A3(new_n407), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n415), .B1(new_n357), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT9), .B(G234), .ZN(new_n427));
  OAI21_X1  g241(.A(G221), .B1(new_n427), .B2(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n368), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G143), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n243), .A2(KEYINPUT82), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n433), .A2(new_n434), .B1(new_n303), .B2(G214), .ZN(new_n435));
  INV_X1    g249(.A(G237), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n218), .A3(G214), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n432), .A2(G143), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT17), .B(G131), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(G214), .A3(new_n303), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT82), .B(G143), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n436), .A2(new_n218), .A3(G214), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(KEYINPUT85), .A3(KEYINPUT17), .A4(G131), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n213), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT86), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n213), .B1(new_n442), .B2(new_n447), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n446), .B(new_n258), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n208), .B(G146), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n446), .A2(new_n459), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n431), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n452), .B2(new_n453), .ZN(new_n465));
  AOI211_X1 g279(.A(KEYINPUT86), .B(new_n213), .C1(new_n442), .C2(new_n447), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n431), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n188), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G475), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n199), .A2(G125), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n204), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT19), .ZN(new_n474));
  AOI21_X1  g288(.A(G146), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n207), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT83), .B(G146), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT84), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n474), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT19), .B1(new_n200), .B2(new_n202), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n211), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n476), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n207), .ZN(new_n486));
  INV_X1    g300(.A(new_n455), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n463), .ZN(new_n489));
  INV_X1    g303(.A(new_n431), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n467), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n470), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G116), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(G116), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n233), .A2(G122), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT89), .B1(new_n505), .B2(KEYINPUT14), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n504), .B(G107), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n501), .A2(new_n505), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n364), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n193), .A2(G143), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT88), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n243), .A2(G128), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n254), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n254), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n507), .B(new_n509), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n512), .B(KEYINPUT13), .Z(new_n517));
  XOR2_X1   g331(.A(new_n510), .B(KEYINPUT88), .Z(new_n518));
  OAI21_X1  g332(.A(G134), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n508), .B(new_n364), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n427), .A2(new_n187), .A3(G953), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n516), .B2(new_n521), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT90), .B(new_n188), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n188), .B1(new_n523), .B2(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT90), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n528), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n431), .B1(new_n488), .B2(new_n463), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n468), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n495), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n494), .B(new_n495), .C1(new_n468), .C2(new_n536), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(KEYINPUT87), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n218), .A2(G952), .ZN(new_n542));
  INV_X1    g356(.A(G234), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n436), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n188), .B(new_n218), .C1(G234), .C2(G237), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n497), .A2(new_n533), .A3(new_n541), .A4(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G210), .B1(G237), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n292), .A2(new_n201), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n201), .B2(new_n284), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n218), .A2(G224), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n557));
  INV_X1    g371(.A(G113), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT5), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n234), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n557), .A2(new_n560), .B1(new_n238), .B2(new_n239), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n375), .B2(new_n376), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n399), .A2(new_n240), .A3(new_n401), .ZN(new_n563));
  XNOR2_X1  g377(.A(G110), .B(G122), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n563), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n564), .B(KEYINPUT78), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n568), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n556), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n252), .A2(G125), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n276), .A2(new_n277), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n278), .A2(new_n283), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n201), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n577));
  INV_X1    g391(.A(new_n555), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n573), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n577), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n553), .B(new_n580), .C1(new_n201), .C2(new_n284), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n565), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n564), .B(KEYINPUT8), .Z(new_n584));
  NAND2_X1  g398(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n238), .A2(new_n586), .A3(KEYINPUT5), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n560), .A2(KEYINPUT80), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n560), .A2(KEYINPUT80), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n238), .A2(new_n239), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n590), .B(new_n591), .C1(new_n375), .C2(new_n376), .ZN(new_n592));
  INV_X1    g406(.A(new_n382), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(new_n561), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n584), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n188), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n552), .B1(new_n572), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n556), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n565), .A2(KEYINPUT6), .B1(new_n567), .B2(new_n568), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n568), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n582), .A2(new_n565), .ZN(new_n602));
  INV_X1    g416(.A(new_n595), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n604), .A3(new_n551), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G214), .B1(G237), .B2(G902), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT77), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n429), .A2(new_n550), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n356), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  NOR2_X1   g427(.A1(new_n429), .A2(new_n232), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n336), .B2(new_n337), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n326), .A2(new_n328), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT91), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT33), .B1(new_n522), .B2(KEYINPUT93), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n523), .B2(new_n524), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n516), .A2(new_n521), .ZN(new_n624));
  INV_X1    g438(.A(new_n522), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n627));
  INV_X1    g441(.A(new_n622), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n526), .A2(G902), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n623), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n623), .A2(new_n629), .A3(new_n631), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT94), .B1(new_n634), .B2(G478), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT95), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n638), .B(new_n632), .C1(new_n633), .C2(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n540), .A2(KEYINPUT87), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n534), .B1(new_n492), .B2(new_n495), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n496), .B(new_n470), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n597), .A2(KEYINPUT92), .A3(new_n605), .ZN(new_n644));
  INV_X1    g458(.A(new_n607), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n551), .B1(new_n601), .B2(new_n604), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT92), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n640), .A2(new_n643), .A3(new_n644), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n548), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND3_X1  g467(.A1(new_n492), .A2(new_n495), .A3(new_n534), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n539), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n470), .A3(new_n532), .A4(new_n549), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT96), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n648), .A2(new_n644), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n539), .A2(new_n654), .B1(G475), .B2(new_n469), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n532), .A4(new_n549), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n657), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n621), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  XNOR2_X1  g481(.A(new_n216), .B(KEYINPUT98), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n229), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n227), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n611), .A2(new_n619), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT37), .B(G110), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n673), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(new_n672), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n341), .B2(new_n355), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n426), .A2(new_n428), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n546), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n544), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n655), .A2(new_n470), .A3(new_n532), .A4(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n658), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n678), .A2(KEYINPUT100), .A3(new_n679), .A4(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n339), .B1(new_n338), .B2(new_n327), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT32), .B(new_n328), .C1(new_n336), .C2(new_n337), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n355), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n679), .A3(new_n672), .A4(new_n684), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  AOI211_X1 g507(.A(KEYINPUT20), .B(new_n538), .C1(new_n491), .C2(new_n467), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n642), .A2(new_n694), .A3(new_n493), .ZN(new_n695));
  INV_X1    g509(.A(G475), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n490), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n698), .B2(new_n467), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n496), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n532), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n645), .A3(new_n672), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT101), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n682), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n679), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n313), .A2(new_n297), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n307), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n334), .A2(new_n335), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n711), .B2(G902), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n686), .B2(new_n687), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n606), .B(KEYINPUT38), .Z(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n703), .A2(new_n707), .A3(new_n708), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  NAND2_X1  g532(.A1(new_n640), .A2(new_n643), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n659), .A4(new_n682), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  INV_X1    g536(.A(new_n682), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n722), .B1(new_n649), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n678), .A2(new_n721), .A3(new_n679), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NAND2_X1  g540(.A1(new_n409), .A2(new_n413), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n188), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n414), .A2(new_n357), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n428), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n356), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n650), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n663), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT104), .B(G116), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G18));
  NOR3_X1   g553(.A1(new_n550), .A2(new_n731), .A3(new_n658), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n688), .A3(new_n672), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n678), .A2(KEYINPUT105), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n323), .A2(new_n324), .A3(new_n301), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n308), .B1(new_n346), .B2(new_n347), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n346), .A2(new_n347), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n336), .B(KEYINPUT106), .C1(new_n751), .C2(new_n308), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n752), .A3(new_n309), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(G472), .C1(new_n326), .C2(G902), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT107), .B1(new_n615), .B2(new_n616), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n327), .A2(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n643), .A2(KEYINPUT108), .A3(new_n532), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT108), .B1(new_n643), .B2(new_n532), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n658), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n731), .A2(new_n548), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n757), .A2(new_n760), .A3(new_n231), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR2_X1   g577(.A1(new_n731), .A2(new_n658), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n719), .A2(new_n723), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n757), .A2(new_n672), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT109), .B(G125), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT42), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n403), .B1(new_n420), .B2(new_n421), .ZN(new_n773));
  INV_X1    g587(.A(new_n408), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n772), .B(new_n406), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n422), .B2(new_n406), .ZN(new_n777));
  OAI211_X1 g591(.A(G469), .B(new_n424), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n415), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n771), .B1(new_n779), .B2(new_n428), .ZN(new_n780));
  INV_X1    g594(.A(new_n428), .ZN(new_n781));
  AOI211_X1 g595(.A(KEYINPUT111), .B(new_n781), .C1(new_n415), .C2(new_n778), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n606), .A2(new_n645), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n688), .A3(new_n231), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n765), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n770), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n688), .A2(new_n231), .A3(new_n784), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n770), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n765), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NOR2_X1   g607(.A1(new_n785), .A2(new_n683), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n254), .ZN(G36));
  INV_X1    g609(.A(new_n643), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n640), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT43), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n672), .B1(new_n617), .B2(new_n618), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n798), .B2(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n784), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n357), .B1(new_n425), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n424), .B1(new_n776), .B2(new_n777), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n806), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n358), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT46), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n730), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n428), .B(new_n705), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n803), .B2(new_n804), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n805), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT114), .B(G137), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G39));
  OAI21_X1  g632(.A(new_n428), .B1(new_n812), .B2(new_n813), .ZN(new_n819));
  AND2_X1   g633(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n822), .B2(new_n820), .ZN(new_n823));
  INV_X1    g637(.A(new_n784), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n786), .A2(new_n688), .A3(new_n231), .A4(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n821), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n199), .ZN(G42));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n658), .B1(new_n701), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n643), .A2(KEYINPUT108), .A3(new_n532), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n682), .B(KEYINPUT119), .Z(new_n832));
  NAND3_X1  g646(.A1(new_n671), .A2(new_n227), .A3(new_n832), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n781), .B(new_n833), .C1(new_n415), .C2(new_n778), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n713), .A2(new_n830), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT120), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n760), .A2(new_n837), .A3(new_n713), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n692), .A2(new_n839), .A3(new_n725), .A4(new_n766), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n725), .A2(new_n766), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n692), .A4(new_n839), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n497), .A2(new_n541), .A3(new_n532), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n606), .A2(new_n549), .A3(new_n609), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT117), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT117), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n614), .A3(new_n619), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n719), .A2(new_n847), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n614), .A2(new_n619), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n612), .A2(new_n850), .A3(new_n673), .A4(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n356), .B(new_n732), .C1(new_n663), .C2(new_n650), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT105), .B1(new_n678), .B2(new_n740), .ZN(new_n855));
  AND4_X1   g669(.A1(KEYINPUT105), .A2(new_n740), .A3(new_n688), .A4(new_n672), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n854), .B(new_n762), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n745), .A2(KEYINPUT116), .A3(new_n762), .A4(new_n854), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n753), .A2(new_n327), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n755), .A2(new_n756), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n672), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n780), .A2(new_n782), .A3(new_n824), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(KEYINPUT118), .A3(new_n765), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n862), .A2(new_n863), .A3(new_n765), .A4(new_n672), .ZN(new_n868));
  INV_X1    g682(.A(new_n780), .ZN(new_n869));
  INV_X1    g683(.A(new_n782), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n784), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n533), .A2(new_n672), .A3(new_n682), .ZN(new_n874));
  INV_X1    g688(.A(new_n660), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n429), .A2(new_n824), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n688), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n785), .B2(new_n683), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n792), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n845), .A2(new_n861), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n842), .B2(new_n844), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n828), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n885), .B2(new_n861), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n878), .B1(new_n791), .B2(new_n787), .ZN(new_n889));
  INV_X1    g703(.A(new_n857), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n853), .A2(new_n883), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n873), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n842), .B2(new_n844), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n888), .A2(new_n893), .A3(KEYINPUT54), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n798), .A2(new_n544), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n231), .A3(new_n757), .ZN(new_n897));
  INV_X1    g711(.A(new_n764), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n542), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n824), .A2(new_n731), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n896), .A2(new_n356), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT48), .Z(new_n902));
  NAND4_X1  g716(.A1(new_n714), .A2(new_n231), .A3(new_n545), .A4(new_n900), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT123), .Z(new_n904));
  AOI211_X1 g718(.A(new_n899), .B(new_n902), .C1(new_n720), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n715), .A2(new_n645), .A3(new_n732), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT50), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT122), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n821), .A2(new_n823), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n729), .A2(new_n730), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n781), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n897), .A2(new_n824), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n896), .A2(new_n864), .A3(new_n900), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n640), .A2(new_n643), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n904), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n910), .A2(new_n916), .A3(KEYINPUT51), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n910), .A2(new_n919), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n913), .B(KEYINPUT121), .Z(new_n922));
  AOI211_X1 g736(.A(new_n824), .B(new_n897), .C1(new_n911), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n905), .B(new_n920), .C1(new_n924), .C2(KEYINPUT51), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n895), .A2(new_n925), .B1(G952), .B2(G953), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n912), .B(KEYINPUT49), .Z(new_n927));
  NAND4_X1  g741(.A1(new_n715), .A2(new_n231), .A3(new_n428), .A4(new_n609), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n927), .A2(new_n928), .A3(new_n797), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n713), .B2(new_n929), .ZN(G75));
  NAND4_X1  g744(.A1(new_n845), .A2(new_n890), .A3(new_n881), .A4(new_n891), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n884), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n599), .A2(new_n600), .A3(new_n598), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n572), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n933), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n218), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n358), .B(KEYINPUT57), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n828), .B1(new_n884), .B2(new_n931), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n894), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n727), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n888), .A2(new_n893), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n188), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n810), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n940), .B1(new_n945), .B2(new_n948), .ZN(G54));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n950));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n932), .A2(G902), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n537), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n940), .B1(new_n952), .B2(new_n537), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n947), .A2(KEYINPUT124), .A3(new_n492), .A4(new_n951), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G60));
  NAND2_X1  g770(.A1(new_n623), .A2(new_n629), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n943), .B2(new_n894), .ZN(new_n961));
  INV_X1    g775(.A(new_n940), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(KEYINPUT125), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  INV_X1    g778(.A(new_n960), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n884), .A2(new_n828), .A3(new_n931), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT54), .B1(new_n888), .B2(new_n893), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n968), .B2(new_n940), .ZN(new_n969));
  INV_X1    g783(.A(new_n959), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n887), .B2(new_n894), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n957), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n963), .A2(new_n969), .A3(new_n972), .ZN(G63));
  INV_X1    g787(.A(new_n224), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n946), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n932), .A2(new_n670), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n979), .A3(new_n962), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G66));
  INV_X1    g796(.A(new_n861), .ZN(new_n983));
  NAND2_X1  g797(.A1(G224), .A2(G953), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n983), .A2(G953), .B1(new_n547), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n570), .B(new_n571), .C1(G898), .C2(new_n218), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(G69));
  AOI21_X1  g801(.A(new_n826), .B1(new_n805), .B2(new_n815), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n356), .A2(new_n760), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n814), .A2(new_n989), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n794), .B(new_n990), .C1(new_n791), .C2(new_n787), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n988), .A2(new_n692), .A3(new_n843), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n473), .A2(new_n474), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n330), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n218), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n843), .A2(new_n717), .A3(new_n692), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT62), .Z(new_n997));
  AOI21_X1  g811(.A(new_n706), .B1(new_n719), .B2(new_n846), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n789), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n1000), .B2(new_n988), .ZN(new_n1001));
  OAI211_X1 g815(.A(G900), .B(new_n995), .C1(new_n1001), .C2(new_n994), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1003), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1005), .B(new_n995), .C1(new_n1001), .C2(new_n994), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(G72));
  XNOR2_X1  g821(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n992), .B2(new_n983), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n307), .A3(new_n300), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n884), .A2(new_n886), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n325), .A2(new_n350), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1013), .A2(new_n1010), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n962), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n349), .A2(new_n308), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n997), .A2(new_n861), .A3(new_n988), .A4(new_n999), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(new_n1010), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1019), .A2(KEYINPUT127), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(KEYINPUT127), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(G57));
endmodule


