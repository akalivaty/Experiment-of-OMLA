//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G197gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT11), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G50gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G43gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT94), .B(KEYINPUT17), .Z(new_n221));
  INV_X1    g020(.A(KEYINPUT93), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n223), .B(new_n224), .C1(new_n222), .C2(new_n216), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(new_n214), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n220), .B(new_n221), .C1(new_n226), .C2(new_n219), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT95), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  AOI21_X1  g029(.A(G1gat), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT96), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n231), .B(new_n233), .Z(new_n234));
  XOR2_X1   g033(.A(KEYINPUT97), .B(G8gat), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n231), .B(new_n233), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT97), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(G8gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n220), .B1(new_n226), .B2(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT98), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n240), .B1(KEYINPUT17), .B2(new_n242), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(new_n228), .B1(new_n246), .B2(new_n240), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT98), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n245), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT99), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT99), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n251), .A2(new_n258), .A3(KEYINPUT18), .A4(new_n245), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n242), .A3(new_n239), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n245), .B(KEYINPUT13), .Z(new_n263));
  AOI21_X1  g062(.A(KEYINPUT100), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  INV_X1    g064(.A(new_n263), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n265), .B(new_n266), .C1(new_n247), .C2(new_n261), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AND4_X1   g068(.A1(new_n208), .A2(new_n255), .A3(new_n260), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n257), .B2(new_n259), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n208), .B1(new_n271), .B2(new_n255), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n260), .A3(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n207), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n208), .A3(new_n255), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(KEYINPUT101), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G228gat), .ZN(new_n279));
  INV_X1    g078(.A(G233gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT81), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G155gat), .B2(G162gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(G155gat), .B2(G162gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT2), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n289), .A3(new_n284), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G197gat), .ZN(new_n306));
  INV_X1    g105(.A(G197gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G204gat), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT75), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT22), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n309), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n304), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n326));
  OAI21_X1  g125(.A(G218gat), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n304), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n329), .A2(KEYINPUT77), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n303), .B1(new_n323), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n329), .B2(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n321), .A2(new_n322), .A3(new_n304), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT78), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n302), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n321), .B2(new_n304), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n304), .B2(new_n321), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n300), .B1(new_n338), .B2(new_n301), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n282), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n298), .A2(new_n289), .A3(new_n284), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n289), .B1(new_n298), .B2(new_n284), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n301), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT78), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT78), .B1(new_n333), .B2(new_n334), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n334), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n301), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n341), .A2(new_n342), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n352), .A3(new_n281), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n340), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT86), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n353), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G22gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n356), .A2(new_n362), .A3(new_n355), .A4(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367));
  OR2_X1    g166(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(G120gat), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT68), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(G120gat), .ZN(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G134gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G127gat), .ZN(new_n378));
  INV_X1    g177(.A(G127gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G134gat), .ZN(new_n380));
  AND2_X1   g179(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n381));
  NOR2_X1   g180(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n378), .B(new_n380), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n372), .A2(G120gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n376), .A2(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n300), .A2(new_n392), .A3(KEYINPUT4), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT71), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n374), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT68), .B1(new_n374), .B2(G113gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n383), .B1(new_n398), .B2(new_n370), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n390), .B1(new_n388), .B2(new_n387), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n381), .A2(new_n382), .ZN(new_n402));
  AND2_X1   g201(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n404), .A3(new_n374), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n373), .A2(new_n375), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n390), .B(new_n402), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n391), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(KEYINPUT71), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n401), .A2(new_n300), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n291), .A2(KEYINPUT3), .A3(new_n299), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n291), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(new_n299), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT83), .B1(new_n399), .B2(new_n400), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n407), .A2(new_n421), .A3(new_n408), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n343), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n413), .B(new_n414), .C1(new_n419), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(G57gat), .B(G85gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n399), .A2(KEYINPUT83), .A3(new_n400), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n421), .B1(new_n407), .B2(new_n408), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n433), .A2(new_n343), .A3(new_n418), .A4(new_n417), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n401), .A2(new_n409), .A3(KEYINPUT4), .A4(new_n300), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n300), .A2(new_n392), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n394), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n434), .A2(new_n414), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n422), .A3(new_n351), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(new_n414), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n413), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n438), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n430), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n429), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n414), .B1(new_n419), .B2(new_n423), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n437), .A2(new_n435), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT84), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n425), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n449), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n367), .B1(new_n448), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n429), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT6), .B1(new_n457), .B2(new_n430), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT85), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n469), .B(KEYINPUT79), .Z(new_n470));
  NAND2_X1  g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471));
  INV_X1    g270(.A(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT66), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G190gat), .ZN(new_n475));
  INV_X1    g274(.A(G183gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT27), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT27), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G183gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n473), .A2(new_n475), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT66), .B(G190gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G183gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(G169gat), .A2(G176gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G169gat), .A2(G176gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n482), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(G169gat), .B2(G176gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n496), .B2(new_n487), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n471), .A2(KEYINPUT24), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(G183gat), .A3(G190gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(G183gat), .A2(G190gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n504), .B2(KEYINPUT65), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n498), .B2(new_n500), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT25), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n484), .A2(new_n476), .B1(new_n498), .B2(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT25), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n497), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n493), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n470), .B1(new_n513), .B2(new_n344), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n482), .A2(new_n486), .A3(new_n492), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n490), .A2(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G169gat), .B2(G176gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n494), .B(new_n517), .C1(new_n506), .C2(new_n507), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n506), .A2(new_n507), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n512), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n470), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n346), .A2(new_n347), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n514), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n332), .A2(new_n335), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n522), .B2(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n470), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n467), .B(new_n468), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n525), .B1(new_n514), .B2(new_n524), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n528), .A2(new_n527), .A3(new_n529), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT80), .B1(new_n539), .B2(KEYINPUT30), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n531), .A2(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n366), .B1(new_n466), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g346(.A1(G227gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT64), .Z(new_n549));
  NOR3_X1   g348(.A1(new_n399), .A2(new_n395), .A3(new_n400), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT71), .B1(new_n407), .B2(new_n408), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n520), .A2(new_n521), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT72), .A4(new_n493), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n401), .A2(new_n409), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n504), .A2(KEYINPUT65), .ZN(new_n556));
  INV_X1    g355(.A(new_n497), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n508), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n512), .B1(new_n558), .B2(new_n511), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n555), .B1(new_n559), .B2(new_n515), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT72), .B1(new_n522), .B2(new_n552), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n549), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(KEYINPUT32), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G15gat), .B(G43gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G99gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n513), .B2(new_n555), .ZN(new_n573));
  INV_X1    g372(.A(new_n549), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n560), .A4(new_n554), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT34), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT32), .B1(new_n569), .B2(new_n564), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n560), .A3(new_n554), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n549), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n554), .A2(new_n560), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n574), .A4(new_n573), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n571), .A2(new_n576), .A3(new_n580), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n583), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n569), .B1(new_n563), .B2(new_n565), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n547), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n584), .C2(new_n587), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(KEYINPUT73), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n585), .B(new_n594), .C1(new_n586), .C2(new_n579), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n593), .A2(KEYINPUT36), .A3(new_n584), .A4(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n546), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n465), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n462), .A2(new_n463), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n459), .A2(KEYINPUT90), .A3(KEYINPUT6), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n534), .B1(new_n531), .B2(KEYINPUT37), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT88), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n537), .A2(new_n538), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g406(.A(KEYINPUT88), .B(KEYINPUT37), .C1(new_n537), .C2(new_n538), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n539), .B1(new_n609), .B2(KEYINPUT38), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT89), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n609), .B2(KEYINPUT38), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n607), .A2(new_n608), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(KEYINPUT89), .A3(new_n614), .A4(new_n603), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n602), .A2(new_n610), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n366), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n414), .B1(new_n411), .B2(new_n434), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT39), .B1(new_n441), .B2(new_n442), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n449), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(KEYINPUT39), .B(new_n414), .C1(new_n411), .C2(new_n434), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n425), .B1(new_n455), .B2(new_n456), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n449), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n627), .B(new_n449), .C1(new_n619), .C2(new_n620), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT87), .B1(new_n628), .B2(new_n618), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT87), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT40), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n625), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n617), .B1(new_n633), .B2(new_n544), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT91), .B1(new_n616), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n465), .A2(new_n598), .B1(new_n462), .B2(new_n463), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n610), .A3(new_n601), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n615), .A2(new_n612), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n634), .B(KEYINPUT91), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n597), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  AND4_X1   g440(.A1(new_n366), .A2(new_n593), .A3(new_n584), .A4(new_n595), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n466), .A3(new_n545), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT35), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT92), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT92), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n646), .A3(KEYINPUT35), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n636), .A2(new_n601), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n544), .A2(new_n588), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n617), .A2(KEYINPUT35), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n278), .B1(new_n641), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G85gat), .A2(G92gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT7), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT8), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n657), .C1(G85gat), .C2(G92gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G99gat), .B(G106gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND3_X1  g459(.A1(new_n228), .A2(new_n243), .A3(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n658), .B(new_n659), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n246), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(G190gat), .B(G218gat), .Z(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT105), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n661), .A2(new_n666), .A3(new_n664), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(G134gat), .B(G162gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT104), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT107), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  INV_X1    g477(.A(new_n670), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n668), .A2(new_n669), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n675), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n679), .A2(new_n680), .B1(new_n666), .B2(new_n665), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n677), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(G71gat), .B(G78gat), .Z(new_n690));
  OR2_X1    g489(.A1(G57gat), .A2(G64gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(G57gat), .A2(G64gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT9), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n699));
  AOI21_X1  g498(.A(G64gat), .B1(KEYINPUT103), .B2(G57gat), .ZN(new_n700));
  OR4_X1    g499(.A1(new_n698), .A2(new_n690), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(KEYINPUT21), .ZN(new_n703));
  NAND2_X1  g502(.A1(G231gat), .A2(G233gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(new_n704), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n379), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n240), .B1(KEYINPUT21), .B2(new_n702), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n705), .B(G127gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n707), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G155gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(G183gat), .B(G211gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n708), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n708), .B2(new_n711), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(G230gat), .A2(G233gat), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n702), .B(new_n663), .C1(new_n721), .C2(new_n659), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT10), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n696), .A2(new_n701), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n659), .A2(new_n721), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n660), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n722), .A2(new_n726), .A3(KEYINPUT109), .A4(new_n723), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n660), .A2(new_n724), .A3(new_n723), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n720), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n726), .ZN(new_n735));
  INV_X1    g534(.A(new_n720), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(G120gat), .B(G148gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(G176gat), .B(G204gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n738), .B(new_n739), .Z(new_n740));
  NAND4_X1  g539(.A1(new_n733), .A2(new_n734), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n742), .B2(new_n736), .ZN(new_n743));
  INV_X1    g542(.A(new_n740), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT110), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n743), .A2(KEYINPUT111), .A3(new_n744), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n743), .B2(new_n744), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n689), .A2(new_n719), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n653), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n466), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n545), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT16), .B(G8gat), .Z(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n760));
  INV_X1    g559(.A(G8gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n756), .ZN(G1325gat));
  OAI21_X1  g561(.A(new_n596), .B1(new_n590), .B2(new_n591), .ZN(new_n763));
  OAI21_X1  g562(.A(G15gat), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n588), .A2(G15gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n753), .B2(new_n765), .ZN(G1326gat));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n366), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT43), .B(G22gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1327gat));
  NAND2_X1  g569(.A1(new_n750), .A2(new_n718), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n689), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n653), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n466), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n209), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT45), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n641), .A2(new_n652), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n677), .A2(new_n683), .A3(new_n687), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n687), .B1(new_n677), .B2(new_n683), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n778), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT44), .B(new_n689), .C1(new_n641), .C2(new_n652), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n275), .A2(new_n276), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT113), .B1(new_n789), .B2(new_n466), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G29gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n789), .A2(KEYINPUT113), .A3(new_n466), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n777), .B1(new_n791), .B2(new_n792), .ZN(G1328gat));
  OAI21_X1  g592(.A(G36gat), .B1(new_n789), .B2(new_n545), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n773), .A2(G36gat), .A3(new_n545), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1329gat));
  OAI21_X1  g596(.A(new_n215), .B1(new_n773), .B2(new_n588), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n592), .A2(G43gat), .A3(new_n596), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g600(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n653), .A2(KEYINPUT114), .A3(new_n772), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n217), .B(new_n617), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n617), .B(new_n788), .C1(new_n783), .C2(new_n784), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G50gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT48), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n804), .B(new_n806), .C1(new_n808), .C2(KEYINPUT48), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1331gat));
  NOR4_X1   g611(.A1(new_n782), .A2(new_n750), .A3(new_n786), .A4(new_n718), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n779), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n775), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g616(.A1(new_n814), .A2(new_n545), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n819));
  AND2_X1   g618(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(G1333gat));
  NOR3_X1   g621(.A1(new_n814), .A2(G71gat), .A3(new_n588), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n814), .A2(new_n763), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(G71gat), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g625(.A1(new_n815), .A2(new_n617), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g627(.A1(new_n787), .A2(new_n718), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n749), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n785), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G85gat), .B1(new_n833), .B2(new_n466), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n643), .A2(new_n646), .A3(KEYINPUT35), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n646), .B1(new_n643), .B2(KEYINPUT35), .ZN(new_n836));
  INV_X1    g635(.A(new_n651), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n600), .A2(new_n367), .B1(KEYINPUT6), .B2(new_n459), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n544), .B1(new_n839), .B2(new_n464), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n763), .B1(new_n840), .B2(new_n366), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT91), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n844), .B2(new_n639), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n831), .B(new_n782), .C1(new_n838), .C2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n750), .A2(G85gat), .A3(new_n466), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n834), .B1(new_n849), .B2(new_n850), .ZN(G1336gat));
  NAND3_X1  g650(.A1(new_n785), .A2(new_n544), .A3(new_n832), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G92gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n750), .A2(G92gat), .A3(new_n545), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n847), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n846), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n852), .A2(G92gat), .B1(new_n860), .B2(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(G1337gat));
  XOR2_X1   g662(.A(KEYINPUT118), .B(G99gat), .Z(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n833), .B2(new_n763), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n750), .A2(new_n588), .A3(new_n864), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n849), .B2(new_n866), .ZN(G1338gat));
  NOR3_X1   g666(.A1(new_n750), .A2(G106gat), .A3(new_n366), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n617), .B(new_n832), .C1(new_n783), .C2(new_n784), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G106gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n859), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n875), .B2(KEYINPUT53), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n877), .B(new_n872), .C1(new_n871), .C2(new_n874), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n873), .B1(new_n876), .B2(new_n878), .ZN(G1339gat));
  NAND2_X1  g678(.A1(new_n742), .A2(new_n736), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n733), .A2(KEYINPUT54), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n742), .A2(new_n736), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n740), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT55), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n746), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n881), .A2(new_n884), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT55), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n890), .B(KEYINPUT55), .C1(new_n881), .C2(new_n884), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n886), .B(new_n786), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n262), .A2(new_n263), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT121), .Z(new_n894));
  NOR2_X1   g693(.A1(new_n251), .A2(new_n245), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n206), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(new_n276), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n749), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n782), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n686), .A2(new_n688), .A3(new_n897), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n886), .B1(new_n889), .B2(new_n891), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n718), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n751), .A2(new_n786), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n617), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n775), .A3(new_n649), .ZN(new_n907));
  OAI21_X1  g706(.A(G113gat), .B1(new_n907), .B2(new_n278), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n903), .A2(new_n905), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(new_n642), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n466), .A2(new_n544), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n786), .A2(new_n368), .A3(new_n369), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(G1340gat));
  OAI21_X1  g713(.A(G120gat), .B1(new_n907), .B2(new_n750), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n749), .A2(new_n374), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n912), .B2(new_n917), .ZN(G1341gat));
  OAI21_X1  g717(.A(G127gat), .B1(new_n907), .B2(new_n718), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n719), .A2(new_n379), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n912), .B2(new_n920), .ZN(G1342gat));
  NAND2_X1  g720(.A1(new_n782), .A2(new_n377), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n912), .A2(KEYINPUT56), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G134gat), .B1(new_n907), .B2(new_n689), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT56), .B1(new_n912), .B2(new_n922), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1343gat));
  NAND2_X1  g725(.A1(new_n887), .A2(new_n888), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n746), .A3(new_n885), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n898), .B1(new_n278), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n689), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n890), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n888), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n782), .A2(new_n933), .A3(new_n897), .A4(new_n886), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n719), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n617), .B1(new_n935), .B2(new_n904), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT57), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n938), .A3(new_n617), .ZN(new_n939));
  INV_X1    g738(.A(new_n278), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n763), .A2(new_n911), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n936), .B2(KEYINPUT57), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n945), .A2(new_n946), .A3(new_n940), .A4(new_n939), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(G141gat), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n366), .B1(new_n903), .B2(new_n905), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(new_n942), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n278), .A2(G141gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT58), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  AND4_X1   g753(.A1(new_n786), .A2(new_n937), .A3(new_n939), .A4(new_n942), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n294), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT58), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n953), .A2(new_n957), .ZN(G1344gat));
  NAND3_X1  g757(.A1(new_n950), .A2(new_n295), .A3(new_n749), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n937), .A2(new_n939), .A3(new_n942), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n295), .C1(new_n960), .C2(new_n749), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n751), .A2(new_n940), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n938), .B(new_n617), .C1(new_n935), .C2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n949), .B2(new_n938), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n942), .A2(new_n749), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n962), .B1(new_n967), .B2(G148gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n959), .B1(new_n961), .B2(new_n968), .ZN(G1345gat));
  AOI21_X1  g768(.A(KEYINPUT124), .B1(new_n950), .B2(new_n719), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(G155gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n950), .A2(KEYINPUT124), .A3(new_n719), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n719), .A2(G155gat), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n971), .A2(new_n972), .B1(new_n960), .B2(new_n973), .ZN(G1346gat));
  INV_X1    g773(.A(G162gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n950), .A2(new_n975), .A3(new_n782), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n960), .A2(new_n782), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n975), .ZN(G1347gat));
  NOR3_X1   g777(.A1(new_n775), .A2(new_n545), .A3(new_n588), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n906), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(G169gat), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n980), .A2(new_n981), .A3(new_n278), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n775), .A2(new_n545), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n910), .A2(new_n786), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n984), .B2(new_n981), .ZN(G1348gat));
  OAI21_X1  g784(.A(G176gat), .B1(new_n980), .B2(new_n750), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n910), .A2(new_n983), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n750), .A2(G176gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(G1349gat));
  NAND4_X1  g788(.A1(new_n910), .A2(new_n485), .A3(new_n719), .A4(new_n983), .ZN(new_n990));
  OAI21_X1  g789(.A(G183gat), .B1(new_n980), .B2(new_n718), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g792(.A1(new_n906), .A2(new_n782), .A3(new_n979), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n994), .A2(new_n995), .A3(G190gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n994), .B2(G190gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n782), .A2(new_n484), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n996), .A2(new_n997), .B1(new_n987), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  OAI221_X1 g800(.A(new_n1001), .B1(new_n987), .B2(new_n998), .C1(new_n996), .C2(new_n997), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1351gat));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n617), .A3(new_n763), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1004), .B1(new_n903), .B2(new_n905), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1005), .A2(new_n307), .A3(new_n786), .ZN(new_n1006));
  XOR2_X1   g805(.A(new_n1006), .B(KEYINPUT126), .Z(new_n1007));
  NAND2_X1  g806(.A1(new_n983), .A2(new_n763), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(new_n940), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n965), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n965), .A2(new_n1011), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1007), .B1(new_n1014), .B2(new_n307), .ZN(G1352gat));
  NAND3_X1  g814(.A1(new_n1005), .A2(new_n305), .A3(new_n749), .ZN(new_n1016));
  XOR2_X1   g815(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  NAND2_X1  g816(.A1(new_n1009), .A2(new_n749), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1018), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1017), .B1(new_n1019), .B2(new_n305), .ZN(G1353gat));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n313), .A3(new_n314), .A4(new_n719), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1008), .A2(new_n718), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g822(.A(G211gat), .B1(new_n965), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g823(.A(KEYINPUT63), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(G1354gat));
  AOI21_X1  g827(.A(G218gat), .B1(new_n1005), .B2(new_n782), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1008), .A2(new_n689), .A3(new_n310), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(G1355gat));
endmodule


