

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n982), .ZN(n850) );
  AND2_X1 U552 ( .A1(n780), .A2(n779), .ZN(n781) );
  BUF_X1 U553 ( .A(n906), .Z(n517) );
  XNOR2_X1 U554 ( .A(n524), .B(n523), .ZN(n906) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NAND2_X1 U556 ( .A1(n906), .A2(G137), .ZN(n525) );
  NAND2_X1 U557 ( .A1(n532), .A2(n531), .ZN(n534) );
  XOR2_X1 U558 ( .A(n739), .B(KEYINPUT31), .Z(n518) );
  XOR2_X1 U559 ( .A(n745), .B(KEYINPUT104), .Z(n519) );
  NOR2_X1 U560 ( .A1(n775), .A2(n774), .ZN(n520) );
  XOR2_X1 U561 ( .A(KEYINPUT29), .B(n727), .Z(n521) );
  XOR2_X1 U562 ( .A(KEYINPUT78), .B(n602), .Z(n522) );
  NAND2_X1 U563 ( .A1(n850), .A2(n712), .ZN(n709) );
  NOR2_X1 U564 ( .A1(n743), .A2(n733), .ZN(n734) );
  BUF_X1 U565 ( .A(n729), .Z(n748) );
  AND2_X1 U566 ( .A1(n747), .A2(n744), .ZN(n745) );
  INV_X1 U567 ( .A(KEYINPUT32), .ZN(n756) );
  XNOR2_X1 U568 ( .A(n757), .B(n756), .ZN(n758) );
  INV_X1 U569 ( .A(KEYINPUT13), .ZN(n591) );
  OR2_X1 U570 ( .A1(n762), .A2(n767), .ZN(n766) );
  XNOR2_X1 U571 ( .A(n591), .B(KEYINPUT74), .ZN(n592) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n796) );
  XNOR2_X1 U573 ( .A(n593), .B(n592), .ZN(n594) );
  INV_X1 U574 ( .A(KEYINPUT17), .ZN(n523) );
  OR2_X1 U575 ( .A1(n821), .A2(n818), .ZN(n837) );
  NOR2_X1 U576 ( .A1(G543), .A2(n556), .ZN(n553) );
  NOR2_X1 U577 ( .A1(G651), .A2(n652), .ZN(n658) );
  NOR2_X2 U578 ( .A1(G543), .A2(G651), .ZN(n664) );
  XNOR2_X1 U579 ( .A(KEYINPUT15), .B(n606), .ZN(n982) );
  AND2_X1 U580 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U581 ( .A(KEYINPUT76), .B(n599), .Z(n976) );
  INV_X1 U582 ( .A(KEYINPUT66), .ZN(n533) );
  NOR2_X1 U583 ( .A1(n541), .A2(n540), .ZN(G164) );
  INV_X1 U584 ( .A(G2105), .ZN(n527) );
  NOR2_X2 U585 ( .A1(G2104), .A2(n527), .ZN(n902) );
  NAND2_X1 U586 ( .A1(n902), .A2(G125), .ZN(n532) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  NAND2_X1 U588 ( .A1(G113), .A2(n901), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n530) );
  AND2_X4 U590 ( .A1(n527), .A2(G2104), .ZN(n905) );
  NAND2_X1 U591 ( .A1(G101), .A2(n905), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT23), .B(n528), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X2 U594 ( .A(n534), .B(n533), .ZN(G160) );
  NAND2_X1 U595 ( .A1(n517), .A2(G138), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G126), .A2(n902), .ZN(n535) );
  XOR2_X1 U597 ( .A(KEYINPUT91), .B(n535), .Z(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G114), .A2(n901), .ZN(n539) );
  NAND2_X1 U600 ( .A1(G102), .A2(n905), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G2446), .B(KEYINPUT106), .ZN(n551) );
  XOR2_X1 U603 ( .A(G2430), .B(G2427), .Z(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT107), .B(G2438), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U606 ( .A(G2435), .B(G2454), .Z(n545) );
  XNOR2_X1 U607 ( .A(G1348), .B(G1341), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U609 ( .A(n547), .B(n546), .Z(n549) );
  XNOR2_X1 U610 ( .A(G2443), .B(G2451), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U613 ( .A1(n552), .A2(G14), .ZN(G401) );
  INV_X1 U614 ( .A(G651), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n553), .Z(n659) );
  NAND2_X1 U616 ( .A1(G64), .A2(n659), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT69), .ZN(n563) );
  XNOR2_X1 U618 ( .A(G543), .B(KEYINPUT0), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT67), .ZN(n652) );
  NOR2_X1 U620 ( .A1(n652), .A2(n556), .ZN(n586) );
  BUF_X1 U621 ( .A(n586), .Z(n663) );
  NAND2_X1 U622 ( .A1(G77), .A2(n663), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G90), .A2(n664), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT9), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G52), .A2(n658), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(G171) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U630 ( .A(G108), .ZN(G238) );
  INV_X1 U631 ( .A(G69), .ZN(G235) );
  NAND2_X1 U632 ( .A1(G75), .A2(n663), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G88), .A2(n664), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G62), .A2(n659), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G50), .A2(n658), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G166) );
  NAND2_X1 U639 ( .A1(n664), .A2(G89), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT4), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G76), .A2(n663), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n573), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G63), .A2(n659), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G51), .A2(n658), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U649 ( .A(n579), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .ZN(n580) );
  XNOR2_X1 U651 ( .A(n580), .B(KEYINPUT79), .ZN(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n581) );
  XOR2_X1 U653 ( .A(n581), .B(KEYINPUT10), .Z(n843) );
  INV_X1 U654 ( .A(n843), .ZN(G223) );
  INV_X1 U655 ( .A(G567), .ZN(n693) );
  NOR2_X1 U656 ( .A1(G223), .A2(n693), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT72), .B(KEYINPUT11), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT71), .B(n584), .Z(G234) );
  NAND2_X1 U660 ( .A1(n659), .A2(G56), .ZN(n585) );
  XNOR2_X1 U661 ( .A(n585), .B(KEYINPUT14), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n586), .A2(G68), .ZN(n587) );
  XNOR2_X1 U663 ( .A(KEYINPUT73), .B(n587), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n664), .A2(G81), .ZN(n588) );
  XOR2_X1 U665 ( .A(n588), .B(KEYINPUT12), .Z(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT75), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G43), .A2(n658), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G860), .A2(n976), .ZN(G153) );
  XNOR2_X1 U672 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n658), .A2(G54), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G79), .A2(n663), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G92), .A2(n664), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n659), .A2(G66), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n522), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U681 ( .A(G868), .ZN(n677) );
  NAND2_X1 U682 ( .A1(n850), .A2(n677), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G65), .A2(n659), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G78), .A2(n663), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G53), .A2(n658), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G91), .A2(n664), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n722) );
  INV_X1 U691 ( .A(n722), .ZN(G299) );
  NOR2_X1 U692 ( .A1(G286), .A2(n677), .ZN(n616) );
  NOR2_X1 U693 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G297) );
  INV_X1 U695 ( .A(G860), .ZN(n634) );
  NAND2_X1 U696 ( .A1(n634), .A2(G559), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n617), .A2(n982), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U699 ( .A1(n982), .A2(G868), .ZN(n619) );
  NOR2_X1 U700 ( .A1(G559), .A2(n619), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n620), .B(KEYINPUT80), .ZN(n622) );
  AND2_X1 U702 ( .A1(n976), .A2(n677), .ZN(n621) );
  NOR2_X1 U703 ( .A1(n622), .A2(n621), .ZN(G282) );
  XOR2_X1 U704 ( .A(G2100), .B(KEYINPUT82), .Z(n632) );
  NAND2_X1 U705 ( .A1(G111), .A2(n901), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G135), .A2(n517), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G123), .A2(n902), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT18), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n626), .B(KEYINPUT81), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n905), .A2(G99), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n935) );
  XOR2_X1 U714 ( .A(G2096), .B(n935), .Z(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U716 ( .A1(G559), .A2(n982), .ZN(n633) );
  XNOR2_X1 U717 ( .A(n633), .B(n976), .ZN(n674) );
  NAND2_X1 U718 ( .A1(n634), .A2(n674), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G67), .A2(n659), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G93), .A2(n664), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G80), .A2(n663), .ZN(n637) );
  XNOR2_X1 U723 ( .A(KEYINPUT83), .B(n637), .ZN(n638) );
  NOR2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n658), .A2(G55), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n676) );
  XNOR2_X1 U727 ( .A(n642), .B(n676), .ZN(G145) );
  NAND2_X1 U728 ( .A1(G73), .A2(n663), .ZN(n643) );
  XNOR2_X1 U729 ( .A(n643), .B(KEYINPUT2), .ZN(n644) );
  XNOR2_X1 U730 ( .A(n644), .B(KEYINPUT84), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G61), .A2(n659), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G48), .A2(n658), .ZN(n648) );
  NAND2_X1 U734 ( .A1(G86), .A2(n664), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U737 ( .A(KEYINPUT85), .B(n651), .ZN(G305) );
  NAND2_X1 U738 ( .A1(G49), .A2(n658), .ZN(n654) );
  NAND2_X1 U739 ( .A1(G87), .A2(n652), .ZN(n653) );
  NAND2_X1 U740 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U741 ( .A1(n659), .A2(n655), .ZN(n657) );
  NAND2_X1 U742 ( .A1(G651), .A2(G74), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(G288) );
  NAND2_X1 U744 ( .A1(n658), .A2(G47), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n659), .A2(G60), .ZN(n660) );
  NAND2_X1 U746 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U747 ( .A(KEYINPUT68), .B(n662), .Z(n668) );
  NAND2_X1 U748 ( .A1(G72), .A2(n663), .ZN(n666) );
  NAND2_X1 U749 ( .A1(G85), .A2(n664), .ZN(n665) );
  AND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(G290) );
  XNOR2_X1 U752 ( .A(KEYINPUT19), .B(G288), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(n676), .ZN(n670) );
  XNOR2_X1 U754 ( .A(G305), .B(n670), .ZN(n672) );
  XOR2_X1 U755 ( .A(G299), .B(G166), .Z(n671) );
  XNOR2_X1 U756 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U757 ( .A(n673), .B(G290), .ZN(n853) );
  XNOR2_X1 U758 ( .A(n674), .B(n853), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n675), .A2(G868), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U762 ( .A(KEYINPUT86), .B(n680), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XNOR2_X1 U764 ( .A(n681), .B(KEYINPUT20), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n682), .B(KEYINPUT87), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n683), .A2(G2090), .ZN(n684) );
  XNOR2_X1 U767 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U769 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U770 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  NAND2_X1 U771 ( .A1(G132), .A2(G82), .ZN(n686) );
  XNOR2_X1 U772 ( .A(n686), .B(KEYINPUT22), .ZN(n687) );
  XNOR2_X1 U773 ( .A(n687), .B(KEYINPUT88), .ZN(n688) );
  NOR2_X1 U774 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U775 ( .A1(G96), .A2(n689), .ZN(n848) );
  NAND2_X1 U776 ( .A1(G2106), .A2(n848), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n690), .B(KEYINPUT89), .ZN(n695) );
  NOR2_X1 U778 ( .A1(G237), .A2(G238), .ZN(n691) );
  NAND2_X1 U779 ( .A1(G120), .A2(n691), .ZN(n692) );
  NOR2_X1 U780 ( .A1(G235), .A2(n692), .ZN(n847) );
  NOR2_X1 U781 ( .A1(n693), .A2(n847), .ZN(n694) );
  NOR2_X1 U782 ( .A1(n695), .A2(n694), .ZN(G319) );
  NAND2_X1 U783 ( .A1(G483), .A2(G661), .ZN(n696) );
  INV_X1 U784 ( .A(G319), .ZN(n919) );
  NOR2_X1 U785 ( .A1(n696), .A2(n919), .ZN(n697) );
  XNOR2_X1 U786 ( .A(n697), .B(KEYINPUT90), .ZN(n846) );
  NAND2_X1 U787 ( .A1(G36), .A2(n846), .ZN(G176) );
  INV_X1 U788 ( .A(G166), .ZN(G303) );
  NAND2_X1 U789 ( .A1(G160), .A2(G40), .ZN(n795) );
  INV_X1 U790 ( .A(n795), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n698), .A2(n796), .ZN(n699) );
  XNOR2_X2 U792 ( .A(n699), .B(KEYINPUT64), .ZN(n729) );
  INV_X1 U793 ( .A(n729), .ZN(n715) );
  XOR2_X1 U794 ( .A(G2078), .B(KEYINPUT101), .Z(n700) );
  XNOR2_X1 U795 ( .A(KEYINPUT25), .B(n700), .ZN(n957) );
  NAND2_X1 U796 ( .A1(n715), .A2(n957), .ZN(n702) );
  INV_X1 U797 ( .A(G1961), .ZN(n981) );
  NAND2_X1 U798 ( .A1(n748), .A2(n981), .ZN(n701) );
  NAND2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n736) );
  NAND2_X1 U800 ( .A1(n736), .A2(G171), .ZN(n728) );
  XNOR2_X1 U801 ( .A(G1996), .B(KEYINPUT103), .ZN(n956) );
  NOR2_X1 U802 ( .A1(n748), .A2(n956), .ZN(n704) );
  XNOR2_X1 U803 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n703) );
  XNOR2_X1 U804 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n748), .A2(G1341), .ZN(n705) );
  NAND2_X1 U806 ( .A1(n706), .A2(n705), .ZN(n711) );
  NAND2_X1 U807 ( .A1(G2067), .A2(n715), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n748), .A2(G1348), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n709), .A2(n976), .ZN(n710) );
  NOR2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U812 ( .A1(n712), .A2(n850), .ZN(n713) );
  NOR2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n721) );
  NAND2_X1 U814 ( .A1(G2072), .A2(n715), .ZN(n716) );
  XNOR2_X1 U815 ( .A(KEYINPUT27), .B(n716), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n729), .A2(G1956), .ZN(n717) );
  XOR2_X1 U817 ( .A(KEYINPUT102), .B(n717), .Z(n718) );
  NOR2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n720) );
  NAND2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n726) );
  OR2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U822 ( .A(n724), .B(KEYINPUT28), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n728), .A2(n521), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n729), .A2(G8), .ZN(n730) );
  XOR2_X1 U826 ( .A(n730), .B(KEYINPUT99), .Z(n774) );
  NOR2_X1 U827 ( .A1(G1966), .A2(n774), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n729), .A2(G2084), .ZN(n731) );
  XNOR2_X1 U829 ( .A(KEYINPUT100), .B(n731), .ZN(n741) );
  INV_X1 U830 ( .A(n741), .ZN(n732) );
  NAND2_X1 U831 ( .A1(n732), .A2(G8), .ZN(n733) );
  XOR2_X1 U832 ( .A(KEYINPUT30), .B(n734), .Z(n735) );
  NOR2_X1 U833 ( .A1(G168), .A2(n735), .ZN(n738) );
  NOR2_X1 U834 ( .A1(G171), .A2(n736), .ZN(n737) );
  NOR2_X1 U835 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U836 ( .A1(n740), .A2(n518), .ZN(n747) );
  AND2_X1 U837 ( .A1(G8), .A2(n741), .ZN(n742) );
  NOR2_X1 U838 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U839 ( .A1(G286), .A2(G8), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n755) );
  INV_X1 U841 ( .A(G8), .ZN(n753) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n774), .ZN(n750) );
  NOR2_X1 U843 ( .A1(n748), .A2(G2090), .ZN(n749) );
  NOR2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n751), .A2(G303), .ZN(n752) );
  OR2_X1 U846 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n519), .A2(n758), .ZN(n773) );
  INV_X1 U849 ( .A(n773), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G166), .A2(G8), .ZN(n759) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  INV_X1 U853 ( .A(n774), .ZN(n767) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n763), .B(KEYINPUT24), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n764), .A2(n767), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n782) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n770) );
  AND2_X1 U859 ( .A1(n770), .A2(KEYINPUT33), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n780) );
  NOR2_X1 U861 ( .A1(G1971), .A2(G303), .ZN(n769) );
  NOR2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n988) );
  INV_X1 U863 ( .A(KEYINPUT33), .ZN(n771) );
  AND2_X1 U864 ( .A1(n988), .A2(n771), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n778) );
  XNOR2_X1 U866 ( .A(G1981), .B(G305), .ZN(n978) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U868 ( .A(n987), .ZN(n775) );
  NOR2_X1 U869 ( .A1(KEYINPUT33), .A2(n520), .ZN(n776) );
  NOR2_X1 U870 ( .A1(n978), .A2(n776), .ZN(n777) );
  AND2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n821) );
  NAND2_X1 U873 ( .A1(G116), .A2(n901), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G128), .A2(n902), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT35), .B(n785), .Z(n792) );
  NAND2_X1 U877 ( .A1(G140), .A2(n517), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n905), .A2(G104), .ZN(n786) );
  XOR2_X1 U879 ( .A(KEYINPUT93), .B(n786), .Z(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT94), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n790), .B(KEYINPUT34), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U884 ( .A(KEYINPUT36), .B(n793), .Z(n915) );
  XOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .Z(n836) );
  NAND2_X1 U886 ( .A1(n915), .A2(n836), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(KEYINPUT95), .ZN(n945) );
  NOR2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n819) );
  NAND2_X1 U889 ( .A1(n945), .A2(n819), .ZN(n826) );
  AND2_X1 U890 ( .A1(KEYINPUT98), .A2(n826), .ZN(n817) );
  NAND2_X1 U891 ( .A1(G107), .A2(n901), .ZN(n798) );
  NAND2_X1 U892 ( .A1(G131), .A2(n517), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G119), .A2(n902), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G95), .A2(n905), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n898) );
  AND2_X1 U898 ( .A1(n898), .A2(G1991), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n902), .A2(G129), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT96), .ZN(n805) );
  NAND2_X1 U901 ( .A1(G117), .A2(n901), .ZN(n804) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U903 ( .A(n806), .B(KEYINPUT97), .ZN(n808) );
  NAND2_X1 U904 ( .A1(G141), .A2(n517), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n905), .A2(G105), .ZN(n809) );
  XOR2_X1 U907 ( .A(KEYINPUT38), .B(n809), .Z(n810) );
  OR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n912) );
  AND2_X1 U909 ( .A1(n912), .A2(G1996), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n822) );
  INV_X1 U911 ( .A(n822), .ZN(n941) );
  XOR2_X1 U912 ( .A(KEYINPUT92), .B(G1986), .Z(n814) );
  XOR2_X1 U913 ( .A(G290), .B(n814), .Z(n995) );
  OR2_X1 U914 ( .A1(n941), .A2(n995), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n815), .A2(n819), .ZN(n816) );
  NAND2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  INV_X1 U917 ( .A(n819), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n837), .A2(n820), .ZN(n841) );
  NOR2_X1 U919 ( .A1(n995), .A2(n821), .ZN(n825) );
  NOR2_X1 U920 ( .A1(KEYINPUT98), .A2(n822), .ZN(n823) );
  AND2_X1 U921 ( .A1(n823), .A2(n826), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n835) );
  INV_X1 U923 ( .A(n826), .ZN(n833) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n912), .ZN(n933) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n827) );
  NOR2_X1 U926 ( .A1(G1991), .A2(n898), .ZN(n937) );
  NOR2_X1 U927 ( .A1(n827), .A2(n937), .ZN(n828) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(n828), .Z(n829) );
  NOR2_X1 U929 ( .A1(n941), .A2(n829), .ZN(n830) );
  NOR2_X1 U930 ( .A1(n933), .A2(n830), .ZN(n831) );
  XOR2_X1 U931 ( .A(KEYINPUT39), .B(n831), .Z(n832) );
  OR2_X1 U932 ( .A1(n833), .A2(n832), .ZN(n834) );
  AND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n839) );
  OR2_X1 U934 ( .A1(n836), .A2(n915), .ZN(n949) );
  AND2_X1 U935 ( .A1(n837), .A2(n949), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U944 ( .A(G132), .ZN(G219) );
  INV_X1 U945 ( .A(G82), .ZN(G220) );
  INV_X1 U946 ( .A(n847), .ZN(n849) );
  NOR2_X1 U947 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U949 ( .A(n976), .B(KEYINPUT114), .ZN(n852) );
  XOR2_X1 U950 ( .A(G171), .B(n850), .Z(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n855) );
  XOR2_X1 U952 ( .A(n853), .B(G286), .Z(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  NOR2_X1 U954 ( .A1(G37), .A2(n856), .ZN(G397) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n859), .B(KEYINPUT111), .Z(n861) );
  XNOR2_X1 U959 ( .A(G1991), .B(G1996), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U961 ( .A(G1976), .B(G1971), .Z(n863) );
  XOR2_X1 U962 ( .A(n981), .B(G1956), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT110), .B(G2474), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(G229) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2678), .B(KEYINPUT43), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT42), .B(G2090), .Z(n871) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2072), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U974 ( .A(G2100), .B(G2096), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n877) );
  XOR2_X1 U976 ( .A(G2078), .B(G2084), .Z(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(G227) );
  NAND2_X1 U978 ( .A1(G124), .A2(n902), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n901), .A2(G112), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G100), .A2(n905), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G136), .A2(n517), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  NAND2_X1 U987 ( .A1(G103), .A2(n905), .ZN(n886) );
  NAND2_X1 U988 ( .A1(G139), .A2(n517), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n901), .A2(G115), .ZN(n887) );
  XNOR2_X1 U991 ( .A(n887), .B(KEYINPUT112), .ZN(n889) );
  NAND2_X1 U992 ( .A1(G127), .A2(n902), .ZN(n888) );
  NAND2_X1 U993 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n926) );
  XNOR2_X1 U996 ( .A(n926), .B(KEYINPUT113), .ZN(n893) );
  XNOR2_X1 U997 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U998 ( .A(G162), .B(G160), .ZN(n895) );
  XNOR2_X1 U999 ( .A(n895), .B(n935), .ZN(n896) );
  XOR2_X1 U1000 ( .A(n897), .B(n896), .Z(n900) );
  XOR2_X1 U1001 ( .A(G164), .B(n898), .Z(n899) );
  XNOR2_X1 U1002 ( .A(n900), .B(n899), .ZN(n917) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n901), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(G130), .A2(n902), .ZN(n903) );
  NAND2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G106), .A2(n905), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(G142), .A2(n517), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1009 ( .A(n909), .B(KEYINPUT45), .Z(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n919), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G397), .A2(n921), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n924), .A2(G395), .ZN(n925) );
  XOR2_X1 U1021 ( .A(n925), .B(KEYINPUT115), .Z(G308) );
  INV_X1 U1022 ( .A(G308), .ZN(G225) );
  INV_X1 U1023 ( .A(G120), .ZN(G236) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1025 ( .A(G2072), .B(n926), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G164), .B(G2078), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(KEYINPUT118), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT119), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n931), .Z(n948) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n934), .Z(n943) );
  XNOR2_X1 U1034 ( .A(G160), .B(G2084), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT116), .B(n939), .Z(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(KEYINPUT117), .B(n946), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n964) );
  XOR2_X1 U1049 ( .A(G2072), .B(G33), .Z(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G28), .ZN(n962) );
  XOR2_X1 U1051 ( .A(n956), .B(G32), .Z(n959) );
  XOR2_X1 U1052 ( .A(n957), .B(G27), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n960), .B(KEYINPUT121), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n965), .B(KEYINPUT53), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(G2090), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G35), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n972), .B(KEYINPUT122), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(G29), .A2(n973), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(KEYINPUT55), .B(n974), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n975), .A2(G11), .ZN(n1030) );
  INV_X1 U1068 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1069 ( .A(n1026), .B(KEYINPUT56), .Z(n1002) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n976), .ZN(n1000) );
  XOR2_X1 U1071 ( .A(G168), .B(G1966), .Z(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT57), .B(n979), .Z(n980) );
  XNOR2_X1 U1074 ( .A(KEYINPUT123), .B(n980), .ZN(n998) );
  XNOR2_X1 U1075 ( .A(G171), .B(n981), .ZN(n984) );
  XOR2_X1 U1076 ( .A(n982), .B(G1348), .Z(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT124), .B(n985), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n991) );
  XOR2_X1 U1081 ( .A(G299), .B(G1956), .Z(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT125), .B(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1028) );
  XOR2_X1 U1090 ( .A(G5), .B(G1961), .Z(n1021) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT126), .B(G4), .Z(n1006) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT60), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(G1986), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(n1014), .B(G24), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(G21), .B(G1966), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

