//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  XOR2_X1   g000(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n187), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n199), .A3(new_n202), .A4(new_n197), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n208), .A3(G143), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n210), .B(G146), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n218), .B(new_n219), .C1(new_n212), .C2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n198), .A2(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n195), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n203), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(G116), .B(G119), .Z(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n230), .A2(new_n232), .B1(KEYINPUT2), .B2(G113), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  INV_X1    g057(.A(new_n240), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n238), .A2(new_n239), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(KEYINPUT67), .A3(new_n240), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n203), .A2(new_n225), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n204), .A2(new_n215), .B1(new_n250), .B2(new_n222), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n248), .B2(new_n251), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n193), .B(new_n242), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n251), .ZN(new_n257));
  INV_X1    g071(.A(new_n241), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n227), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT65), .B1(new_n251), .B2(KEYINPUT30), .ZN(new_n261));
  AND4_X1   g075(.A1(KEYINPUT65), .A2(new_n216), .A3(KEYINPUT30), .A4(new_n226), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT66), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n216), .A2(KEYINPUT65), .A3(KEYINPUT30), .A4(new_n226), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT66), .B1(new_n269), .B2(new_n260), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n257), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n193), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n256), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT70), .B(G902), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n227), .A2(new_n247), .A3(new_n246), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n252), .B2(new_n253), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G472), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(G472), .C1(new_n273), .C2(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n257), .A2(new_n193), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n286), .B1(new_n289), .B2(new_n263), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n292), .A2(new_n293), .B1(new_n241), .B2(new_n227), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n290), .A2(new_n291), .B1(new_n193), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n291), .B(new_n296), .C1(new_n264), .C2(new_n270), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n285), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n294), .A2(new_n193), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n296), .B1(new_n264), .B2(new_n270), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(KEYINPUT31), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n297), .A2(new_n298), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT69), .B1(new_n290), .B2(new_n291), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n284), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n275), .B2(G234), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(G119), .B(G128), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT72), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT24), .B(G110), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G119), .B2(new_n217), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT23), .A3(G128), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n321), .A2(new_n323), .B1(G119), .B2(new_n217), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n317), .A2(new_n319), .B1(G110), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n327));
  AND2_X1   g141(.A1(G125), .A2(G140), .ZN(new_n328));
  NOR2_X1   g142(.A1(G125), .A2(G140), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n208), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT16), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n332), .A2(KEYINPUT16), .A3(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n333), .A3(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n326), .A2(new_n327), .A3(new_n330), .A4(new_n336), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n317), .A2(new_n319), .B1(G110), .B2(new_n324), .ZN(new_n338));
  AOI21_X1  g152(.A(G146), .B1(new_n331), .B2(new_n333), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT22), .B(G137), .Z(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT75), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n346), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n337), .B2(new_n341), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n315), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT76), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT25), .B1(new_n352), .B2(new_n274), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n275), .C1(new_n347), .C2(new_n349), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n314), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT9), .B(G234), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G221), .B1(new_n360), .B2(G902), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT77), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n213), .A2(new_n214), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n364), .B2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G104), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(G107), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n365), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT79), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n368), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(G101), .A3(new_n373), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n363), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n204), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n367), .A2(G104), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n364), .A2(G107), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n371), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT10), .A3(new_n222), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n222), .A2(new_n371), .A3(new_n384), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n380), .A2(new_n381), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n189), .A2(G227), .ZN(new_n392));
  INV_X1    g206(.A(G140), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G110), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n394), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G110), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT10), .B1(new_n386), .B2(new_n222), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n379), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n381), .B1(new_n404), .B2(new_n387), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT80), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n219), .A2(new_n218), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n212), .A2(new_n221), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n385), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n388), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(KEYINPUT12), .A3(new_n204), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n411), .B2(new_n204), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND4_X1   g228(.A1(KEYINPUT10), .A2(new_n222), .A3(new_n371), .A4(new_n384), .ZN(new_n415));
  NOR4_X1   g229(.A1(new_n379), .A2(new_n403), .A3(new_n415), .A4(new_n204), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n407), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n385), .B(new_n222), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n381), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(KEYINPUT12), .A3(new_n204), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n401), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n406), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G469), .B1(new_n426), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n402), .A2(new_n414), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n375), .A2(G101), .A3(new_n373), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n376), .B2(new_n374), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n387), .B(new_n390), .C1(new_n431), .C2(new_n363), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n204), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n401), .B1(new_n433), .B2(new_n391), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n428), .B(new_n275), .C1(new_n429), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n425), .B1(new_n405), .B2(new_n416), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n422), .A2(new_n401), .A3(new_n391), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n274), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n362), .B1(new_n427), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT82), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n377), .A2(new_n378), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n241), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n322), .A3(G116), .ZN(new_n452));
  OAI211_X1 g266(.A(G113), .B(new_n452), .C1(new_n236), .C2(new_n451), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n386), .A2(new_n240), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n448), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n377), .A2(new_n378), .B1(new_n237), .B2(new_n240), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n240), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n385), .ZN(new_n458));
  INV_X1    g272(.A(new_n446), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT6), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n447), .B1(new_n456), .B2(new_n458), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n215), .A2(G125), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n222), .A2(new_n332), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n189), .A2(G224), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n457), .A2(new_n472), .A3(new_n385), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n457), .B2(new_n385), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n454), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n446), .B(KEYINPUT8), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT7), .B(new_n469), .C1(new_n468), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT84), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT84), .B1(new_n466), .B2(new_n467), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n480), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n486));
  INV_X1    g300(.A(new_n477), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n457), .A2(new_n385), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n473), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n490), .B2(new_n454), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(new_n480), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n460), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n471), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n471), .A2(new_n495), .A3(new_n497), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n445), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT91), .B1(new_n217), .B2(G143), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n210), .A3(G128), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(new_n504), .B1(new_n217), .B2(G143), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n195), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  INV_X1    g321(.A(G116), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(G122), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT90), .A3(G116), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n367), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(G107), .A3(new_n513), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(KEYINPUT14), .A3(G107), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n514), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n502), .A2(new_n504), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n217), .A2(G143), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n195), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n505), .A2(G134), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n526), .A3(G134), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n512), .A2(G107), .A3(new_n513), .ZN(new_n529));
  AOI21_X1  g343(.A(G107), .B1(new_n512), .B2(new_n513), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n521), .A2(new_n526), .A3(G134), .A4(new_n522), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n520), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n360), .A2(new_n313), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n520), .B2(new_n533), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n520), .A2(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT92), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n275), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G478), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI221_X1 g361(.A(new_n275), .B1(KEYINPUT15), .B2(new_n545), .C1(new_n540), .C2(new_n543), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n332), .A2(new_n393), .ZN(new_n551));
  NAND2_X1  g365(.A1(G125), .A2(G140), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(G146), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n330), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(KEYINPUT18), .A2(G131), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G143), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(G143), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G214), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n562), .A2(G237), .A3(G953), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n210), .A2(KEYINPUT86), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n556), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n210), .A2(KEYINPUT86), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n556), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n558), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n555), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G131), .B1(new_n561), .B2(new_n565), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n202), .A3(new_n570), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n328), .B2(new_n329), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n551), .A2(KEYINPUT19), .A3(new_n552), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n573), .A2(new_n574), .B1(new_n579), .B2(new_n208), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n572), .B1(new_n580), .B2(new_n336), .ZN(new_n581));
  XNOR2_X1  g395(.A(G113), .B(G122), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n364), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n550), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n566), .A2(new_n571), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n554), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n561), .A2(new_n565), .A3(G131), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n202), .B1(new_n568), .B2(new_n570), .ZN(new_n588));
  OAI22_X1  g402(.A1(new_n587), .A2(new_n588), .B1(new_n578), .B2(G146), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n334), .B(KEYINPUT74), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n583), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT87), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n573), .A2(new_n574), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n340), .A2(new_n339), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n583), .A3(new_n586), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n584), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G475), .ZN(new_n601));
  INV_X1    g415(.A(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n598), .A2(new_n586), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n592), .A2(KEYINPUT88), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n592), .A4(new_n586), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT89), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT89), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n602), .A4(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G475), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n600), .A2(KEYINPUT20), .A3(new_n601), .A4(new_n602), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n189), .A2(G952), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(G234), .B2(G237), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n189), .B(new_n275), .C1(G234), .C2(G237), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT21), .B(G898), .Z(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n549), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n443), .A2(new_n501), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n312), .A2(new_n358), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT93), .B(G101), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G3));
  NAND2_X1  g443(.A1(new_n299), .A2(new_n300), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n303), .B1(new_n630), .B2(new_n307), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n310), .A2(new_n275), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(G472), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n471), .A2(new_n495), .A3(new_n497), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n497), .B1(new_n471), .B2(new_n495), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n444), .B(new_n623), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n540), .B2(new_n543), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n538), .B1(new_n536), .B2(new_n539), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n542), .A2(new_n537), .A3(new_n535), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(KEYINPUT33), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(G478), .A3(new_n275), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n544), .A2(new_n545), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n616), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n636), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n633), .A2(new_n358), .A3(new_n646), .A4(new_n443), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(new_n616), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n549), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n633), .A2(new_n358), .A3(new_n652), .A4(new_n443), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n342), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n315), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n356), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n626), .A2(new_n633), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT37), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n399), .ZN(G12));
  INV_X1    g476(.A(new_n659), .ZN(new_n663));
  AOI211_X1 g477(.A(new_n285), .B(new_n303), .C1(new_n630), .C2(new_n307), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT32), .B1(new_n310), .B2(new_n302), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n666), .B2(new_n284), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n443), .A2(new_n501), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n618), .B1(new_n620), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT94), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT94), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n667), .A2(new_n674), .A3(new_n668), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n670), .B(KEYINPUT39), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n362), .B(new_n678), .C1(new_n427), .C2(new_n442), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT40), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n193), .B1(new_n276), .B2(new_n257), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n602), .B1(new_n290), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G472), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n659), .B1(new_n666), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n634), .A2(new_n635), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT38), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n549), .A2(new_n616), .A3(new_n444), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n680), .A2(new_n684), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR2_X1   g504(.A1(new_n645), .A2(new_n670), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n667), .A2(new_n668), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  OR2_X1    g507(.A1(new_n439), .A2(new_n428), .ZN(new_n694));
  INV_X1    g508(.A(new_n362), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n440), .B1(new_n439), .B2(new_n428), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT95), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n439), .A2(new_n428), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n436), .B2(new_n441), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT95), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n695), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n312), .A2(new_n704), .A3(new_n358), .A4(new_n646), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n312), .A2(new_n704), .A3(new_n358), .A4(new_n652), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n703), .A3(new_n501), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT96), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n699), .A2(new_n703), .A3(KEYINPUT96), .A4(new_n501), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n667), .A3(new_n625), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XOR2_X1   g531(.A(KEYINPUT98), .B(G472), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n306), .A2(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n277), .A2(new_n272), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n630), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n632), .A2(new_n718), .B1(new_n302), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n685), .A2(new_n687), .A3(new_n624), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n704), .A2(new_n358), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  AND2_X1   g539(.A1(new_n714), .A2(new_n691), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n722), .A2(new_n659), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n311), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n631), .A2(KEYINPUT100), .A3(KEYINPUT32), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n284), .A3(new_n733), .A4(new_n304), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n358), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT99), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n696), .A2(new_n697), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n422), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT80), .B1(new_n422), .B2(new_n391), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n425), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n406), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n428), .B1(new_n742), .B2(new_n602), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n736), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n427), .A2(new_n442), .A3(KEYINPUT99), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n362), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n499), .A2(new_n444), .A3(new_n500), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n645), .A3(new_n670), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n748), .A3(KEYINPUT42), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n730), .B1(new_n735), .B2(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n746), .A2(new_n748), .A3(KEYINPUT42), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT101), .A3(new_n358), .A4(new_n734), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n357), .B1(new_n666), .B2(new_n284), .ZN(new_n753));
  INV_X1    g567(.A(new_n747), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n691), .A3(new_n754), .A4(new_n746), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n750), .A2(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT102), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  AND4_X1   g573(.A1(new_n312), .A2(new_n746), .A3(new_n358), .A4(new_n754), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT103), .B1(new_n760), .B2(new_n671), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n312), .A2(new_n746), .A3(new_n358), .A4(new_n754), .ZN(new_n762));
  INV_X1    g576(.A(new_n671), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n195), .ZN(G36));
  NAND2_X1  g581(.A1(new_n426), .A2(KEYINPUT45), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT104), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n769), .B(G469), .C1(KEYINPUT45), .C2(new_n426), .ZN(new_n770));
  NAND2_X1  g584(.A1(G469), .A2(G902), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n737), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n771), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n362), .B(new_n678), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n650), .A2(new_n644), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n633), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n659), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n747), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n776), .B(new_n784), .C1(new_n783), .C2(new_n782), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  AOI21_X1  g600(.A(new_n362), .B1(new_n774), .B2(new_n775), .ZN(new_n787));
  NAND2_X1  g601(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n312), .A2(new_n358), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(new_n791), .A3(new_n748), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  INV_X1    g608(.A(new_n704), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n747), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n619), .B1(new_n779), .B2(new_n780), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n727), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n722), .A2(new_n358), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n686), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n445), .A3(new_n803), .A4(new_n704), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n789), .A2(new_n791), .B1(new_n362), .B2(new_n701), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(new_n754), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT112), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n799), .B(new_n806), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n796), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n666), .A2(new_n683), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n812), .A2(new_n813), .A3(new_n357), .A4(new_n619), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n650), .A3(new_n643), .A4(new_n642), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n804), .A2(new_n816), .A3(KEYINPUT50), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n807), .A2(new_n809), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n820), .B2(KEYINPUT114), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n811), .A3(new_n815), .A4(new_n817), .ZN(new_n824));
  INV_X1    g638(.A(new_n735), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n798), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  AOI21_X1  g641(.A(new_n617), .B1(new_n827), .B2(KEYINPUT48), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n645), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n814), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n801), .B1(new_n712), .B2(new_n713), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  INV_X1    g650(.A(new_n670), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT108), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n687), .B(new_n685), .C1(KEYINPUT108), .C2(new_n837), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n684), .A2(new_n746), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n676), .A2(new_n728), .A3(new_n692), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n673), .A2(new_n675), .B1(new_n726), .B2(new_n727), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n692), .A4(new_n840), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n549), .A2(new_n616), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n312), .A2(new_n443), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n746), .A2(new_n722), .A3(new_n830), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n663), .B(new_n747), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n760), .A2(KEYINPUT103), .A3(new_n671), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n764), .B1(new_n762), .B2(new_n763), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n850), .A2(new_n837), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n750), .A2(new_n752), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n755), .A2(new_n756), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n715), .A2(new_n705), .A3(new_n708), .A4(new_n724), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n660), .A2(new_n653), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n627), .A2(new_n647), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT106), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n627), .A2(new_n862), .A3(new_n647), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n853), .A2(new_n856), .A3(new_n858), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT107), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n859), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n627), .A2(new_n862), .A3(new_n647), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n862), .B1(new_n627), .B2(new_n647), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n857), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(KEYINPUT107), .A3(new_n856), .A4(new_n853), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n869), .A2(new_n875), .B1(new_n843), .B2(new_n845), .ZN(new_n876));
  XNOR2_X1  g690(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n836), .B(new_n867), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT109), .B1(new_n876), .B2(KEYINPUT53), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n757), .A2(new_n873), .A3(new_n857), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT107), .B1(new_n881), .B2(new_n853), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n861), .A2(new_n863), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n705), .A2(new_n708), .A3(new_n724), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n715), .A3(new_n884), .A4(new_n870), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n848), .A2(new_n849), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n659), .A3(new_n837), .A4(new_n754), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n761), .B2(new_n765), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n885), .A2(new_n888), .A3(new_n757), .A4(new_n868), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n846), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT109), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n876), .A2(new_n877), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n880), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI211_X1 g709(.A(KEYINPUT111), .B(new_n879), .C1(KEYINPUT54), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n898), .B2(new_n878), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n833), .B(new_n835), .C1(new_n896), .C2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(G952), .A2(G953), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n701), .B(KEYINPUT49), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n803), .A2(new_n358), .A3(new_n778), .A4(new_n903), .ZN(new_n904));
  OR4_X1    g718(.A1(new_n362), .A2(new_n904), .A3(new_n445), .A4(new_n813), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(G75));
  NAND2_X1  g720(.A1(new_n869), .A2(new_n875), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n877), .B1(new_n907), .B2(new_n846), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n867), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n274), .A3(new_n498), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n465), .B(new_n470), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  NOR2_X1   g727(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n914));
  AND2_X1   g728(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n911), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n189), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n913), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(KEYINPUT116), .B(new_n913), .C1(new_n911), .C2(new_n919), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n916), .B(new_n918), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(G51));
  INV_X1    g739(.A(new_n867), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n908), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n928), .A3(new_n878), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n908), .C2(new_n926), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n771), .B(KEYINPUT57), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n930), .A4(new_n931), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n934), .B(new_n935), .C1(new_n434), .C2(new_n429), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n910), .A2(new_n274), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(new_n770), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n917), .B1(new_n936), .B2(new_n938), .ZN(G54));
  NAND4_X1  g753(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .A4(new_n274), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n600), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n917), .ZN(G60));
  AND2_X1   g756(.A1(new_n638), .A2(new_n641), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n896), .A2(new_n899), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n943), .A2(new_n947), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n929), .A2(new_n930), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n918), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(KEYINPUT120), .A3(new_n918), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n948), .A2(new_n955), .ZN(G63));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n909), .B2(new_n867), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n657), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n918), .ZN(new_n962));
  INV_X1    g776(.A(new_n352), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  INV_X1    g780(.A(new_n964), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n917), .B1(new_n960), .B2(new_n657), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n957), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT121), .B1(new_n962), .B2(new_n964), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n966), .A3(new_n968), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(G66));
  NAND2_X1  g788(.A1(new_n885), .A2(new_n189), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n622), .A2(G224), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(KEYINPUT122), .B2(new_n975), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n461), .B(new_n464), .C1(G898), .C2(new_n189), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G69));
  OAI21_X1  g796(.A(new_n269), .B1(KEYINPUT30), .B2(new_n251), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n578), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n793), .A2(new_n785), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n685), .A2(new_n687), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n776), .A2(new_n986), .A3(new_n825), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n676), .A2(new_n728), .A3(new_n692), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n856), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n989), .A2(new_n766), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(G953), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n189), .A2(G900), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n990), .A2(new_n689), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n651), .A2(new_n645), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n753), .A2(new_n679), .A3(new_n754), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n998), .A2(new_n985), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n189), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n995), .B1(new_n984), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT123), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n1001), .B2(new_n885), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n271), .B(KEYINPUT125), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1009), .A2(new_n193), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT126), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n992), .A2(new_n874), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1008), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n272), .B(new_n1010), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n271), .A2(new_n272), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n895), .B(new_n1008), .C1(new_n290), .C2(new_n1018), .ZN(new_n1019));
  AND4_X1   g833(.A1(new_n918), .A2(new_n1013), .A3(new_n1016), .A4(new_n1019), .ZN(G57));
endmodule


