

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G1966), .A2(n788), .ZN(n683) );
  NAND2_X1 U549 ( .A1(n515), .A2(n753), .ZN(n792) );
  NOR2_X1 U550 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U551 ( .A1(n722), .A2(G1341), .ZN(n513) );
  NAND2_X1 U552 ( .A1(n785), .A2(n808), .ZN(n514) );
  XOR2_X1 U553 ( .A(n752), .B(KEYINPUT101), .Z(n515) );
  AND2_X1 U554 ( .A1(n737), .A2(n685), .ZN(n686) );
  BUF_X1 U555 ( .A(n689), .Z(n722) );
  INV_X1 U556 ( .A(KEYINPUT96), .ZN(n682) );
  NAND2_X1 U557 ( .A1(n680), .A2(n783), .ZN(n681) );
  XNOR2_X1 U558 ( .A(n681), .B(KEYINPUT64), .ZN(n689) );
  NAND2_X1 U559 ( .A1(n689), .A2(G8), .ZN(n788) );
  INV_X1 U560 ( .A(n1014), .ZN(n753) );
  INV_X1 U561 ( .A(G2104), .ZN(n521) );
  NOR2_X1 U562 ( .A1(n514), .A2(n790), .ZN(n791) );
  NAND2_X1 U563 ( .A1(n516), .A2(G2104), .ZN(n517) );
  NAND2_X1 U564 ( .A1(n792), .A2(n791), .ZN(n815) );
  NOR2_X1 U565 ( .A1(G651), .A2(n622), .ZN(n647) );
  INV_X1 U566 ( .A(G2105), .ZN(n516) );
  XNOR2_X2 U567 ( .A(n517), .B(KEYINPUT67), .ZN(n869) );
  NAND2_X1 U568 ( .A1(G102), .A2(n869), .ZN(n520) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n518), .Z(n597) );
  NAND2_X1 U571 ( .A1(G138), .A2(n597), .ZN(n519) );
  NAND2_X1 U572 ( .A1(n520), .A2(n519), .ZN(n526) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NAND2_X1 U574 ( .A1(G114), .A2(n874), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n521), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U576 ( .A(n522), .B(KEYINPUT65), .ZN(n875) );
  NAND2_X1 U577 ( .A1(G126), .A2(n875), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U580 ( .A1(n869), .A2(G101), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(KEYINPUT68), .Z(n527) );
  XNOR2_X1 U582 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G125), .A2(n875), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n529), .B(KEYINPUT66), .ZN(n530) );
  AND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n679) );
  NAND2_X1 U586 ( .A1(G137), .A2(n597), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G113), .A2(n874), .ZN(n532) );
  AND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n677) );
  AND2_X1 U589 ( .A1(n679), .A2(n677), .ZN(G160) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U591 ( .A(G57), .ZN(G237) );
  INV_X1 U592 ( .A(G132), .ZN(G219) );
  INV_X1 U593 ( .A(G82), .ZN(G220) );
  INV_X1 U594 ( .A(G651), .ZN(n538) );
  NOR2_X1 U595 ( .A1(G543), .A2(n538), .ZN(n534) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n534), .Z(n640) );
  NAND2_X1 U597 ( .A1(G64), .A2(n640), .ZN(n536) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NAND2_X1 U599 ( .A1(G52), .A2(n647), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT70), .B(n537), .ZN(n543) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U603 ( .A1(G90), .A2(n639), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n622), .A2(n538), .ZN(n643) );
  NAND2_X1 U605 ( .A1(G77), .A2(n643), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(G171) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  NAND2_X1 U610 ( .A1(G89), .A2(n639), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT4), .B(n544), .Z(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT75), .ZN(n547) );
  NAND2_X1 U613 ( .A1(G76), .A2(n643), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G63), .A2(n640), .ZN(n550) );
  NAND2_X1 U617 ( .A1(G51), .A2(n647), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n557) );
  INV_X1 U626 ( .A(G223), .ZN(n822) );
  NAND2_X1 U627 ( .A1(G567), .A2(n822), .ZN(n556) );
  XNOR2_X1 U628 ( .A(n557), .B(n556), .ZN(G234) );
  NAND2_X1 U629 ( .A1(n640), .A2(G56), .ZN(n558) );
  XOR2_X1 U630 ( .A(KEYINPUT14), .B(n558), .Z(n565) );
  NAND2_X1 U631 ( .A1(n639), .A2(G81), .ZN(n559) );
  XNOR2_X1 U632 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U633 ( .A1(G68), .A2(n643), .ZN(n560) );
  NAND2_X1 U634 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(n562), .ZN(n563) );
  XNOR2_X1 U636 ( .A(KEYINPUT73), .B(n563), .ZN(n564) );
  NOR2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n647), .A2(G43), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n998) );
  INV_X1 U640 ( .A(G860), .ZN(n589) );
  OR2_X1 U641 ( .A1(n998), .A2(n589), .ZN(G153) );
  INV_X1 U642 ( .A(G868), .ZN(n658) );
  NOR2_X1 U643 ( .A1(G301), .A2(n658), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G92), .A2(n639), .ZN(n569) );
  NAND2_X1 U645 ( .A1(G79), .A2(n643), .ZN(n568) );
  NAND2_X1 U646 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U647 ( .A1(G66), .A2(n640), .ZN(n571) );
  NAND2_X1 U648 ( .A1(G54), .A2(n647), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U651 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n574) );
  XNOR2_X1 U652 ( .A(n575), .B(n574), .ZN(n892) );
  NOR2_X1 U653 ( .A1(n892), .A2(G868), .ZN(n576) );
  NOR2_X1 U654 ( .A1(n577), .A2(n576), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G65), .A2(n640), .ZN(n579) );
  NAND2_X1 U656 ( .A1(G53), .A2(n647), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G91), .A2(n639), .ZN(n581) );
  NAND2_X1 U659 ( .A1(G78), .A2(n643), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n584), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U663 ( .A(KEYINPUT76), .B(n658), .ZN(n585) );
  NOR2_X1 U664 ( .A1(G286), .A2(n585), .ZN(n588) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n586) );
  XOR2_X1 U666 ( .A(KEYINPUT77), .B(n586), .Z(n587) );
  NOR2_X1 U667 ( .A1(n588), .A2(n587), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n589), .A2(G559), .ZN(n590) );
  INV_X1 U669 ( .A(n892), .ZN(n995) );
  NAND2_X1 U670 ( .A1(n590), .A2(n995), .ZN(n591) );
  XNOR2_X1 U671 ( .A(n591), .B(KEYINPUT78), .ZN(n592) );
  XNOR2_X1 U672 ( .A(KEYINPUT16), .B(n592), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n998), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n995), .A2(G868), .ZN(n593) );
  NOR2_X1 U675 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G123), .A2(n875), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT18), .ZN(n600) );
  BUF_X1 U679 ( .A(n597), .Z(n870) );
  NAND2_X1 U680 ( .A1(G135), .A2(n870), .ZN(n598) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(n598), .Z(n599) );
  NAND2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G99), .A2(n869), .ZN(n602) );
  NAND2_X1 U684 ( .A1(G111), .A2(n874), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n966) );
  XNOR2_X1 U687 ( .A(n966), .B(G2096), .ZN(n606) );
  INV_X1 U688 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(G156) );
  XNOR2_X1 U690 ( .A(n998), .B(KEYINPUT80), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n995), .A2(G559), .ZN(n607) );
  XNOR2_X1 U692 ( .A(n608), .B(n607), .ZN(n656) );
  NOR2_X1 U693 ( .A1(G860), .A2(n656), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G93), .A2(n639), .ZN(n610) );
  NAND2_X1 U695 ( .A1(G80), .A2(n643), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U697 ( .A(n611), .B(KEYINPUT81), .ZN(n613) );
  NAND2_X1 U698 ( .A1(G55), .A2(n647), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n640), .A2(G67), .ZN(n614) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n614), .Z(n615) );
  OR2_X1 U702 ( .A1(n616), .A2(n615), .ZN(n659) );
  XOR2_X1 U703 ( .A(n617), .B(n659), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n647), .ZN(n619) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U707 ( .A1(n640), .A2(n620), .ZN(n621) );
  XOR2_X1 U708 ( .A(KEYINPUT83), .B(n621), .Z(n624) );
  NAND2_X1 U709 ( .A1(n622), .A2(G87), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G88), .A2(n639), .ZN(n626) );
  NAND2_X1 U712 ( .A1(G75), .A2(n643), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n640), .A2(G62), .ZN(n627) );
  XOR2_X1 U715 ( .A(KEYINPUT84), .B(n627), .Z(n628) );
  NOR2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n647), .A2(G50), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G72), .A2(n643), .ZN(n633) );
  NAND2_X1 U721 ( .A1(G60), .A2(n640), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G85), .A2(n639), .ZN(n634) );
  XNOR2_X1 U724 ( .A(KEYINPUT69), .B(n634), .ZN(n635) );
  NOR2_X1 U725 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n647), .A2(G47), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U728 ( .A1(G86), .A2(n639), .ZN(n642) );
  NAND2_X1 U729 ( .A1(G61), .A2(n640), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U732 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n647), .A2(G48), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(G305) );
  XOR2_X1 U736 ( .A(n659), .B(G288), .Z(n654) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(G299), .ZN(n650) );
  XNOR2_X1 U738 ( .A(n650), .B(G290), .ZN(n651) );
  XNOR2_X1 U739 ( .A(G166), .B(n651), .ZN(n652) );
  XNOR2_X1 U740 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n654), .B(n653), .ZN(n889) );
  XNOR2_X1 U742 ( .A(KEYINPUT85), .B(n889), .ZN(n655) );
  XNOR2_X1 U743 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X1 U744 ( .A1(n658), .A2(n657), .ZN(n661) );
  NOR2_X1 U745 ( .A1(G868), .A2(n659), .ZN(n660) );
  NOR2_X1 U746 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n666) );
  XNOR2_X1 U754 ( .A(KEYINPUT22), .B(n666), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n667), .A2(G96), .ZN(n668) );
  NOR2_X1 U756 ( .A1(G218), .A2(n668), .ZN(n669) );
  XOR2_X1 U757 ( .A(KEYINPUT86), .B(n669), .Z(n828) );
  NAND2_X1 U758 ( .A1(n828), .A2(G2106), .ZN(n673) );
  NAND2_X1 U759 ( .A1(G120), .A2(G108), .ZN(n670) );
  NOR2_X1 U760 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U761 ( .A1(G69), .A2(n671), .ZN(n827) );
  NAND2_X1 U762 ( .A1(G567), .A2(n827), .ZN(n672) );
  NAND2_X1 U763 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U764 ( .A(KEYINPUT87), .B(n674), .ZN(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n826) );
  NAND2_X1 U768 ( .A1(n826), .A2(G36), .ZN(G176) );
  AND2_X1 U769 ( .A1(n677), .A2(G40), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n782) );
  INV_X1 U771 ( .A(n782), .ZN(n680) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n783) );
  XNOR2_X1 U773 ( .A(n683), .B(n682), .ZN(n737) );
  INV_X1 U774 ( .A(G8), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n722), .A2(G2084), .ZN(n735) );
  NOR2_X1 U776 ( .A1(n684), .A2(n735), .ZN(n685) );
  XOR2_X1 U777 ( .A(KEYINPUT30), .B(n686), .Z(n687) );
  NOR2_X1 U778 ( .A1(G168), .A2(n687), .ZN(n688) );
  XNOR2_X1 U779 ( .A(n688), .B(KEYINPUT99), .ZN(n693) );
  XOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .Z(n942) );
  NOR2_X1 U781 ( .A1(n722), .A2(n942), .ZN(n691) );
  INV_X1 U782 ( .A(n689), .ZN(n704) );
  NOR2_X1 U783 ( .A1(G1961), .A2(n704), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n695), .A2(G301), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U788 ( .A1(n695), .A2(G301), .ZN(n696) );
  XNOR2_X1 U789 ( .A(KEYINPUT97), .B(n696), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n704), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U791 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n697) );
  XNOR2_X1 U792 ( .A(n698), .B(n697), .ZN(n700) );
  INV_X1 U793 ( .A(G1956), .ZN(n917) );
  NOR2_X1 U794 ( .A1(n704), .A2(n917), .ZN(n699) );
  NOR2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n715) );
  INV_X1 U796 ( .A(G299), .ZN(n714) );
  NAND2_X1 U797 ( .A1(n715), .A2(n714), .ZN(n713) );
  NAND2_X1 U798 ( .A1(n704), .A2(G1996), .ZN(n701) );
  XNOR2_X1 U799 ( .A(n701), .B(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n998), .A2(n513), .ZN(n702) );
  AND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n709), .A2(n995), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n722), .A2(G1348), .ZN(n706) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n704), .ZN(n705) );
  NAND2_X1 U805 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n711) );
  AND2_X1 U807 ( .A1(n995), .A2(n709), .ZN(n710) );
  NOR2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n718) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U811 ( .A(n716), .B(KEYINPUT28), .Z(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U813 ( .A(KEYINPUT29), .B(n719), .Z(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n733) );
  NOR2_X1 U815 ( .A1(n722), .A2(G2090), .ZN(n724) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n788), .ZN(n723) );
  NOR2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n725), .A2(G303), .ZN(n727) );
  AND2_X1 U819 ( .A1(n733), .A2(n727), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n734), .A2(n726), .ZN(n731) );
  INV_X1 U821 ( .A(n727), .ZN(n728) );
  OR2_X1 U822 ( .A1(n728), .A2(G286), .ZN(n729) );
  AND2_X1 U823 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n732), .B(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G8), .A2(n735), .ZN(n736) );
  AND2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n755) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  AND2_X1 U831 ( .A1(n755), .A2(n1004), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n754), .A2(n740), .ZN(n745) );
  INV_X1 U833 ( .A(n1004), .ZN(n743) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n1007), .A2(n741), .ZN(n742) );
  OR2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U839 ( .A1(n746), .A2(n788), .ZN(n747) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n747), .ZN(n748) );
  XNOR2_X1 U841 ( .A(n748), .B(KEYINPUT100), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n1007), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U843 ( .A1(n788), .A2(n749), .ZN(n750) );
  XNOR2_X1 U844 ( .A(G1981), .B(G305), .ZN(n1014) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n758) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U847 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n788), .A2(n759), .ZN(n785) );
  NAND2_X1 U850 ( .A1(G141), .A2(n870), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G117), .A2(n874), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n869), .A2(G105), .ZN(n762) );
  XNOR2_X1 U854 ( .A(n762), .B(KEYINPUT38), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G129), .A2(n875), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  OR2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n882) );
  NOR2_X1 U858 ( .A1(G1996), .A2(n882), .ZN(n974) );
  NAND2_X1 U859 ( .A1(G107), .A2(n874), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G119), .A2(n875), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U862 ( .A(KEYINPUT94), .B(n769), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G95), .A2(n869), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G131), .A2(n870), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n862) );
  INV_X1 U867 ( .A(G1991), .ZN(n939) );
  NOR2_X1 U868 ( .A1(n862), .A2(n939), .ZN(n775) );
  AND2_X1 U869 ( .A1(n882), .A2(G1996), .ZN(n774) );
  NOR2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n978) );
  INV_X1 U871 ( .A(n978), .ZN(n779) );
  NOR2_X1 U872 ( .A1(G1986), .A2(G290), .ZN(n776) );
  AND2_X1 U873 ( .A1(n939), .A2(n862), .ZN(n967) );
  NOR2_X1 U874 ( .A1(n776), .A2(n967), .ZN(n777) );
  XNOR2_X1 U875 ( .A(n777), .B(KEYINPUT102), .ZN(n778) );
  NOR2_X1 U876 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U877 ( .A1(n974), .A2(n780), .ZN(n781) );
  XNOR2_X1 U878 ( .A(KEYINPUT39), .B(n781), .ZN(n784) );
  NOR2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n817) );
  NAND2_X1 U880 ( .A1(n784), .A2(n817), .ZN(n808) );
  NOR2_X1 U881 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XNOR2_X1 U882 ( .A(n786), .B(KEYINPUT24), .ZN(n787) );
  XNOR2_X1 U883 ( .A(n787), .B(KEYINPUT95), .ZN(n789) );
  NOR2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .Z(n816) );
  XNOR2_X1 U886 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n807) );
  NAND2_X1 U887 ( .A1(n870), .A2(G140), .ZN(n793) );
  XNOR2_X1 U888 ( .A(KEYINPUT89), .B(n793), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n869), .A2(G104), .ZN(n794) );
  XOR2_X1 U890 ( .A(n794), .B(KEYINPUT88), .Z(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U892 ( .A(KEYINPUT90), .B(n797), .Z(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT34), .B(n798), .Z(n805) );
  NAND2_X1 U894 ( .A1(G128), .A2(n875), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n874), .A2(G116), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT91), .B(n799), .Z(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U898 ( .A(n802), .B(KEYINPUT92), .ZN(n803) );
  XNOR2_X1 U899 ( .A(KEYINPUT35), .B(n803), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U901 ( .A(n807), .B(n806), .Z(n886) );
  AND2_X1 U902 ( .A1(n816), .A2(n886), .ZN(n984) );
  NAND2_X1 U903 ( .A1(n984), .A2(n817), .ZN(n813) );
  INV_X1 U904 ( .A(n808), .ZN(n811) );
  XOR2_X1 U905 ( .A(G1986), .B(G290), .Z(n996) );
  NAND2_X1 U906 ( .A1(n978), .A2(n996), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n809), .A2(n817), .ZN(n810) );
  OR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n816), .A2(n886), .ZN(n980) );
  NAND2_X1 U912 ( .A1(n980), .A2(n817), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  XOR2_X1 U914 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n820) );
  XNOR2_X1 U915 ( .A(n821), .B(n820), .ZN(G329) );
  NAND2_X1 U916 ( .A1(n822), .A2(G2106), .ZN(n823) );
  XOR2_X1 U917 ( .A(KEYINPUT105), .B(n823), .Z(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U919 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G108), .B(KEYINPUT111), .ZN(G238) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  NOR2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(G2100), .B(G2096), .Z(n830) );
  XNOR2_X1 U929 ( .A(KEYINPUT42), .B(G2678), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2090), .Z(n832) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1986), .B(G1976), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1961), .B(G1971), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n839), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(G2474), .B(G1981), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1956), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(G229) );
  NAND2_X1 U947 ( .A1(G136), .A2(n870), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G112), .A2(n874), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G124), .A2(n875), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n869), .A2(G100), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U954 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U955 ( .A1(G118), .A2(n874), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G130), .A2(n875), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n870), .A2(G142), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n855), .B(KEYINPUT106), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G106), .A2(n869), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U962 ( .A(KEYINPUT107), .B(n858), .ZN(n859) );
  XNOR2_X1 U963 ( .A(KEYINPUT45), .B(n859), .ZN(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n866) );
  XOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n864) );
  XNOR2_X1 U966 ( .A(G164), .B(n862), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U969 ( .A(G160), .B(n966), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G103), .A2(n869), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT108), .B(n873), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G115), .A2(n874), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G127), .A2(n875), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n962) );
  XOR2_X1 U980 ( .A(n881), .B(n962), .Z(n884) );
  XOR2_X1 U981 ( .A(n882), .B(G162), .Z(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U984 ( .A1(G37), .A2(n887), .ZN(n888) );
  XOR2_X1 U985 ( .A(KEYINPUT109), .B(n888), .Z(G395) );
  XNOR2_X1 U986 ( .A(G286), .B(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n998), .B(G171), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n894) );
  XOR2_X1 U989 ( .A(n892), .B(KEYINPUT110), .Z(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U992 ( .A(KEYINPUT104), .B(G2446), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2454), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n898), .B(G2451), .Z(n900) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2435), .B(G2427), .Z(n902) );
  XNOR2_X1 U999 ( .A(G2430), .B(G2438), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(G1348), .B(KEYINPUT59), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n912), .B(G4), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G19), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(G1981), .B(G6), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n920) );
  XOR2_X1 U1018 ( .A(G20), .B(n917), .Z(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT126), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT60), .B(n921), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G21), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G5), .B(G1961), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G22), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(G23), .B(G1976), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n929) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(KEYINPUT58), .B(n930), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n933) );
  XNOR2_X1 U1034 ( .A(n934), .B(n933), .ZN(n936) );
  INV_X1 U1035 ( .A(G16), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1037 ( .A1(n937), .A2(G11), .ZN(n994) );
  XNOR2_X1 U1038 ( .A(KEYINPUT119), .B(G2090), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(G35), .ZN(n954) );
  XOR2_X1 U1040 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n952) );
  XOR2_X1 U1041 ( .A(G2072), .B(G33), .Z(n941) );
  XNOR2_X1 U1042 ( .A(n939), .B(G25), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1046 ( .A(G32), .B(G1996), .Z(n945) );
  NAND2_X1 U1047 ( .A1(n945), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(G2067), .ZN(n946) );
  XNOR2_X1 U1049 ( .A(G26), .B(n946), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n952), .B(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G34), .B(G2084), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(KEYINPUT122), .B(n958), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(n960), .B(KEYINPUT55), .ZN(n992) );
  XNOR2_X1 U1060 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G164), .B(G2078), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(n961), .B(KEYINPUT117), .ZN(n964) );
  XOR2_X1 U1063 ( .A(G2072), .B(n962), .Z(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(KEYINPUT50), .B(n965), .ZN(n987) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT112), .B(n968), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(G160), .B(G2084), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1070 ( .A(KEYINPUT113), .B(n971), .ZN(n982) );
  XOR2_X1 U1071 ( .A(G2090), .B(G162), .Z(n972) );
  XNOR2_X1 U1072 ( .A(KEYINPUT114), .B(n972), .ZN(n973) );
  NOR2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n975) );
  XNOR2_X1 U1075 ( .A(n976), .B(n975), .ZN(n977) );
  NAND2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT116), .B(n985), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n989), .B(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(G29), .A2(n990), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1022) );
  XNOR2_X1 U1086 ( .A(KEYINPUT56), .B(G16), .ZN(n1019) );
  XNOR2_X1 U1087 ( .A(G1348), .B(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1012) );
  XNOR2_X1 U1089 ( .A(n998), .B(G1341), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G301), .B(G1961), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G166), .B(G1971), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT123), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(KEYINPUT124), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(G168), .B(G1966), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT125), .B(n1020), .Z(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

