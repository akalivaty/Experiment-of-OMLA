//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(G2105), .B2(new_n473), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n476), .A2(G124), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n463), .A2(new_n465), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n475), .A2(KEYINPUT69), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n480), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(new_n482), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n482), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT70), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n475), .A2(new_n495), .A3(G126), .A4(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT4), .B1(new_n483), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n475), .A2(new_n500), .A3(G138), .A4(new_n482), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OR3_X1    g084(.A1(new_n508), .A2(KEYINPUT71), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n508), .B2(new_n509), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT72), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n514), .B(new_n516), .C1(new_n505), .C2(new_n506), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(new_n521), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND2_X1   g101(.A1(new_n507), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT74), .B(G89), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n514), .A2(new_n516), .A3(G64), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(G52), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n522), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(new_n541), .C1(new_n522), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n540), .B1(new_n544), .B2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n537), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n508), .A2(new_n550), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT78), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT77), .B(KEYINPUT8), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT79), .Z(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n508), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n507), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n523), .A2(G91), .ZN(new_n569));
  INV_X1    g144(.A(G78), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n570), .A2(new_n513), .A3(KEYINPUT80), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT80), .B1(new_n570), .B2(new_n513), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n514), .A2(new_n516), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n568), .A2(new_n569), .A3(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n544), .A2(new_n546), .ZN(new_n578));
  INV_X1    g153(.A(new_n540), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT81), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  AOI211_X1 g156(.A(new_n581), .B(new_n540), .C1(new_n544), .C2(new_n546), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G301));
  NAND2_X1  g159(.A1(new_n527), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G87), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n527), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n523), .A2(G86), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n537), .C2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n523), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n527), .A2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G60), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n574), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT82), .B1(new_n597), .B2(G651), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n593), .B(new_n594), .C1(new_n600), .C2(new_n601), .ZN(G290));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OR3_X1    g178(.A1(new_n522), .A2(KEYINPUT84), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT84), .B1(new_n522), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n537), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n527), .A2(G54), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n608), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n583), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT83), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(KEYINPUT83), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(KEYINPUT83), .B2(new_n617), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n568), .A2(new_n569), .A3(new_n576), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n614), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g204(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  INV_X1    g206(.A(new_n487), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G135), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n633), .A2(KEYINPUT87), .B1(G123), .B2(new_n476), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n482), .B2(G111), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n634), .B1(KEYINPUT87), .B2(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n483), .A2(new_n462), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  NAND2_X1  g215(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n638), .B(new_n643), .C1(KEYINPUT86), .C2(G2100), .ZN(G156));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT88), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n651), .B(new_n656), .Z(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT89), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT17), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n665), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT90), .Z(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n669), .A2(new_n663), .A3(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT91), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT92), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT93), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(KEYINPUT94), .A3(new_n680), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n679), .A2(new_n680), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n685), .A3(new_n681), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n686), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n690), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT95), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G23), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT33), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1976), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(G6), .ZN(new_n711));
  INV_X1    g286(.A(G305), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT96), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n705), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n705), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT97), .B(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n710), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n705), .A2(G24), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G290), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n632), .A2(G131), .ZN(new_n729));
  OR2_X1    g304(.A1(G95), .A2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G107), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n462), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n476), .A2(G119), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n725), .B2(new_n724), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n721), .B2(KEYINPUT34), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n722), .A2(new_n726), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n637), .A2(new_n727), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT102), .Z(new_n745));
  NAND2_X1  g320(.A1(G168), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G16), .B2(G21), .ZN(new_n747));
  INV_X1    g322(.A(G1966), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(new_n752), .B(G160), .S(G29), .Z(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n553), .B2(G16), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G1341), .ZN(new_n758));
  INV_X1    g333(.A(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT30), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT30), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n760), .A2(new_n761), .A3(new_n727), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n749), .A2(new_n755), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n747), .A2(new_n748), .B1(G1341), .B2(new_n757), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n753), .A2(new_n754), .ZN(new_n765));
  NOR2_X1   g340(.A1(G5), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G171), .B2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G1961), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n727), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n727), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n705), .A2(G20), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT23), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT23), .B1(new_n622), .B2(new_n705), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n774), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  NOR4_X1   g356(.A1(new_n763), .A2(new_n773), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n727), .A2(G26), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(G116), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n462), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n476), .A2(G128), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n485), .A2(new_n486), .A3(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n727), .ZN(new_n791));
  MUX2_X1   g366(.A(new_n783), .B(new_n791), .S(KEYINPUT28), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT99), .B(G2067), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G32), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n632), .A2(G141), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NOR2_X1   g373(.A1(new_n462), .A2(G2105), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n476), .A2(G129), .B1(G105), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n796), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT27), .B(G1996), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n614), .B2(G16), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT98), .B(G1348), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1961), .ZN(new_n810));
  INV_X1    g385(.A(new_n767), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n782), .A2(new_n794), .A3(new_n805), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n485), .A2(new_n486), .A3(G139), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT100), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n485), .A2(new_n486), .A3(new_n816), .A4(G139), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n799), .A2(G103), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT25), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n815), .A2(KEYINPUT101), .A3(new_n819), .A4(new_n817), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n475), .A2(G127), .ZN(new_n825));
  NAND2_X1  g400(.A1(G115), .A2(G2104), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n482), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  MUX2_X1   g404(.A(G33), .B(new_n829), .S(G29), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2072), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n727), .A2(G35), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G162), .B2(new_n727), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT29), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(G2090), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT103), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n834), .A2(G2090), .B1(new_n778), .B2(new_n779), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n813), .A2(new_n831), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n743), .A2(new_n745), .A3(new_n839), .ZN(G311));
  NAND3_X1  g415(.A1(new_n743), .A2(new_n745), .A3(new_n839), .ZN(G150));
  AOI22_X1  g416(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n537), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n508), .A2(new_n845), .B1(new_n846), .B2(new_n522), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n613), .A2(new_n625), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT104), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n843), .B2(new_n847), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n553), .A3(new_n857), .ZN(new_n858));
  OAI221_X1 g433(.A(new_n856), .B1(new_n549), .B2(new_n552), .C1(new_n843), .C2(new_n847), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n854), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n861), .B2(G860), .ZN(G145));
  NAND2_X1  g437(.A1(new_n476), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(new_n482), .B2(G118), .ZN(new_n865));
  INV_X1    g440(.A(G142), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n863), .B1(new_n864), .B2(new_n865), .C1(new_n487), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n640), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n734), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n829), .A2(new_n790), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n824), .A2(new_n828), .A3(new_n789), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n801), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n789), .B1(new_n824), .B2(new_n828), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n827), .B(new_n790), .C1(new_n822), .C2(new_n823), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n802), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n873), .A2(new_n876), .A3(G164), .ZN(new_n877));
  AOI21_X1  g452(.A(G164), .B1(new_n873), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n503), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n873), .A2(new_n876), .A3(G164), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n869), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n488), .B(G160), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n637), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n869), .A2(KEYINPUT107), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n877), .B2(new_n878), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n881), .A2(new_n882), .A3(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(new_n887), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n888), .A2(new_n894), .A3(KEYINPUT108), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(G395));
  XNOR2_X1  g479(.A(new_n598), .B(new_n599), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(G288), .A3(new_n593), .A4(new_n594), .ZN(new_n906));
  NAND2_X1  g481(.A1(G290), .A2(new_n707), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(new_n907), .A3(G303), .ZN(new_n908));
  AOI21_X1  g483(.A(G303), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(G305), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G166), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n907), .A3(G303), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n712), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT109), .Z(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT110), .Z(new_n919));
  AND2_X1   g494(.A1(new_n858), .A2(new_n859), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n627), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n611), .A2(new_n612), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n622), .A2(new_n922), .A3(new_n610), .A4(new_n608), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n613), .A2(G299), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT41), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n923), .B2(new_n924), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n921), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n917), .A2(new_n919), .A3(new_n927), .A4(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n919), .A2(new_n917), .B1(new_n927), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n849), .A2(new_n616), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  OAI21_X1  g513(.A(G168), .B1(new_n580), .B2(new_n582), .ZN(new_n939));
  NAND2_X1  g514(.A1(G286), .A2(G171), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(G286), .A2(G171), .A3(KEYINPUT112), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n920), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n860), .A2(new_n942), .A3(new_n939), .A4(new_n943), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(KEYINPUT113), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n920), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n930), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT114), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n945), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n926), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n947), .A2(new_n930), .A3(new_n954), .A4(new_n949), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n951), .A2(new_n915), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n910), .A2(new_n914), .A3(KEYINPUT115), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT115), .B1(new_n910), .B2(new_n914), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n931), .A2(new_n952), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n925), .B1(new_n947), .B2(new_n949), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n962), .A3(new_n895), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n959), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n895), .A3(new_n956), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n964), .B(KEYINPUT44), .C1(new_n967), .C2(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n956), .A2(new_n962), .A3(new_n969), .A4(new_n895), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n503), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n469), .B(KEYINPUT68), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n980));
  OAI21_X1  g555(.A(G2105), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n466), .A2(new_n467), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n482), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(G40), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(G160), .A2(KEYINPUT116), .A3(G40), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n978), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n789), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n802), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT127), .Z(new_n994));
  NOR2_X1   g569(.A1(new_n990), .A2(G1996), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n990), .A2(G1986), .A3(G290), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n801), .B(G1996), .Z(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n992), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n735), .A2(new_n738), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n734), .A2(new_n737), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n989), .B2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n1002), .A2(new_n1004), .B1(G2067), .B2(new_n789), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n989), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  NOR3_X1   g585(.A1(new_n998), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n984), .B(KEYINPUT116), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n591), .B2(new_n537), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G1981), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n591), .A2(new_n537), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n589), .A3(new_n1019), .A4(new_n590), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G305), .A2(G1981), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1021), .A3(KEYINPUT49), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1015), .B(new_n1024), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G288), .A2(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1014), .A2(new_n1032), .A3(G8), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1015), .A2(new_n1032), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1029), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G303), .A2(G8), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1039), .B(KEYINPUT55), .Z(new_n1040));
  NOR2_X1   g615(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n977), .B(G1384), .C1(new_n497), .C2(new_n502), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n988), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(G1971), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n986), .B(new_n987), .C1(new_n1013), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1013), .A2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1047), .A2(KEYINPUT117), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1044), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1038), .A2(G8), .A3(new_n1040), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n707), .A2(new_n1030), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT121), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1029), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1015), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(G8), .A3(new_n1040), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1038), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1012), .A2(new_n754), .A3(new_n1063), .A4(new_n1049), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(G168), .C1(new_n1043), .C2(G1966), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G168), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1040), .B1(new_n1054), .B2(G8), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1062), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1055), .B(new_n1060), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1071), .A3(G168), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1012), .A2(new_n978), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n748), .ZN(new_n1076));
  AOI21_X1  g651(.A(G168), .B1(new_n1076), .B2(new_n1064), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  OAI211_X1 g653(.A(G8), .B(new_n1065), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1012), .A2(new_n771), .A3(new_n978), .A4(new_n1074), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n810), .B1(new_n1046), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT53), .A3(new_n771), .A4(new_n1012), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1079), .A2(new_n1091), .A3(new_n1080), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1082), .A2(new_n583), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1046), .B2(new_n1086), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1012), .A2(new_n991), .A3(new_n1013), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n613), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT124), .B(G2072), .Z(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT56), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1043), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1012), .A2(KEYINPUT122), .A3(new_n1063), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1046), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1086), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1104), .B2(G1956), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G299), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1097), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1100), .B(new_n1107), .C1(new_n1104), .C2(G1956), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1095), .A2(new_n613), .A3(new_n1096), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1097), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1095), .A2(new_n1096), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1110), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1104), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n779), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1100), .A4(new_n1107), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1014), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(new_n1125), .B1(new_n1075), .B2(G1996), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n553), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT59), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1112), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n984), .A2(new_n1084), .A3(G2078), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1088), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1085), .A2(new_n1087), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1130), .A2(G301), .B1(new_n1133), .B2(G171), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1134), .A2(KEYINPUT54), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1090), .A2(new_n583), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1085), .A2(new_n1132), .A3(G301), .A4(new_n1087), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT125), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1141), .B(KEYINPUT54), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1073), .B(new_n1093), .C1(new_n1129), .C2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1044), .B1(new_n1120), .B2(G2090), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1040), .B1(new_n1145), .B2(G8), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1062), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1072), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1006), .ZN(new_n1149));
  XNOR2_X1  g724(.A(G290), .B(new_n725), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n990), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1011), .B1(new_n1148), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g727(.A1(G227), .A2(new_n460), .ZN(new_n1154));
  AND2_X1   g728(.A1(new_n965), .A2(new_n959), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n956), .A2(new_n895), .ZN(new_n1156));
  OAI21_X1  g730(.A(KEYINPUT43), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1157), .B2(new_n970), .ZN(new_n1158));
  OAI21_X1  g732(.A(new_n703), .B1(new_n658), .B2(new_n657), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n1159), .B1(new_n898), .B2(new_n899), .ZN(new_n1160));
  AND2_X1   g734(.A1(new_n1158), .A2(new_n1160), .ZN(G308));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(G225));
endmodule


