//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OAI21_X1  g0006(.A(new_n205), .B1(new_n206), .B2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G13), .ZN(new_n208));
  NAND4_X1  g0008(.A1(new_n208), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G250), .B1(G257), .B2(G264), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G68), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n206), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n221), .B(new_n234), .C1(KEYINPUT0), .C2(new_n213), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G97), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n253), .A2(KEYINPUT66), .B1(G77), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(G1698), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT67), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(KEYINPUT66), .B2(new_n253), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(G226), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n214), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n269), .B2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n284), .A2(new_n286), .B1(new_n201), .B2(new_n215), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n215), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT8), .B(G58), .Z(new_n291));
  AOI21_X1  g0091(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n279), .A2(new_n214), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n282), .B1(G50), .B2(new_n283), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n268), .A2(new_n295), .A3(new_n275), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n278), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n268), .A2(G190), .A3(new_n275), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n294), .B(KEYINPUT9), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(G200), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n288), .B(KEYINPUT68), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n202), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n285), .A2(G50), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(G20), .B2(new_n230), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n310), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n280), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OR3_X1    g0115(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n317));
  AOI22_X1  g0117(.A1(G68), .A2(new_n281), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n313), .B2(new_n314), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n229), .A2(G1698), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n251), .B(new_n321), .C1(G226), .C2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n267), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(new_n272), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n273), .B2(new_n231), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n266), .B1(new_n322), .B2(new_n323), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT13), .B1(new_n331), .B2(new_n328), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(G179), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT71), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n325), .B2(new_n329), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n331), .A2(new_n328), .A3(KEYINPUT13), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(G169), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n320), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G200), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n330), .B2(new_n332), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT69), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(G190), .A3(new_n332), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n315), .A2(new_n319), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(KEYINPUT69), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n327), .B1(new_n273), .B2(new_n223), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n258), .A2(new_n229), .A3(G1698), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G107), .B2(new_n258), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n261), .B2(new_n231), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n354), .B2(new_n267), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n281), .A2(G77), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G77), .B2(new_n283), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n291), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT15), .B(G87), .Z(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n215), .A3(G33), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n293), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n355), .B2(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n355), .A2(new_n295), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT67), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n260), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G238), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n266), .B1(new_n371), .B2(new_n353), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n277), .B1(new_n372), .B2(new_n351), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n368), .A2(new_n373), .A3(new_n365), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AND4_X1   g0175(.A1(new_n306), .A2(new_n350), .A3(new_n367), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n251), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G68), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n228), .A2(new_n230), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n218), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n285), .A2(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n230), .B1(new_n378), .B2(new_n379), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n385), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(new_n280), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n291), .A2(new_n283), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n281), .B2(new_n291), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n255), .A2(new_n257), .A3(G223), .A4(new_n252), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT72), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n251), .A2(new_n397), .A3(G223), .A4(new_n252), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n251), .A2(G226), .A3(G1698), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n396), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n267), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n272), .B1(new_n274), .B2(G232), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G190), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(KEYINPUT73), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n408), .A3(new_n267), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n394), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT17), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n394), .B(new_n413), .C1(new_n404), .C2(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n391), .A2(new_n393), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n403), .A2(new_n295), .ZN(new_n417));
  INV_X1    g0217(.A(new_n409), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n408), .B1(new_n401), .B2(new_n267), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n402), .A2(new_n403), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n277), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n416), .A2(new_n420), .A3(KEYINPUT18), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n422), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(new_n394), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n407), .A2(new_n409), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n417), .B1(new_n277), .B2(new_n421), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n430), .A2(KEYINPUT74), .A3(KEYINPUT18), .A4(new_n416), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n415), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n376), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT6), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n438), .A2(new_n224), .A3(G107), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n438), .B2(new_n248), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n440), .A2(new_n215), .B1(new_n202), .B2(new_n286), .ZN(new_n441));
  INV_X1    g0241(.A(G107), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n378), .B2(new_n379), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n280), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n283), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n269), .A2(G33), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n293), .A2(new_n283), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(G97), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n255), .A2(new_n257), .A3(G250), .A4(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n251), .A2(KEYINPUT77), .A3(G250), .A4(G1698), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT4), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n251), .A2(G244), .A3(new_n252), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n451), .A2(new_n452), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n455), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(new_n252), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n267), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n269), .A2(G45), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n266), .B(G257), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT79), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n466), .A2(new_n468), .B1(new_n264), .B2(new_n265), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n264), .A2(new_n265), .B1(new_n269), .B2(G45), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT79), .B(G257), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n470), .A2(new_n271), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(new_n466), .A3(new_n468), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n464), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n444), .B(new_n448), .C1(new_n480), .C2(new_n405), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n267), .C1(new_n458), .C2(new_n463), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n482), .B1(new_n487), .B2(new_n343), .ZN(new_n488));
  INV_X1    g0288(.A(new_n486), .ZN(new_n489));
  AND4_X1   g0289(.A1(G244), .A2(new_n255), .A3(new_n257), .A4(new_n252), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n455), .B1(new_n450), .B2(new_n449), .ZN(new_n491));
  INV_X1    g0291(.A(new_n457), .ZN(new_n492));
  AND4_X1   g0292(.A1(G250), .A2(new_n255), .A3(new_n257), .A4(G1698), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(KEYINPUT77), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n494), .A3(new_n462), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n485), .B1(new_n495), .B2(new_n267), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n295), .B(new_n479), .C1(new_n489), .C2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n480), .A2(new_n277), .B1(new_n444), .B2(new_n448), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n488), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n283), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n293), .A2(new_n283), .A3(new_n446), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n457), .B(new_n215), .C1(G33), .C2(new_n224), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(G20), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n280), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  OAI221_X1 g0313(.A(new_n505), .B1(new_n504), .B2(new_n506), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n266), .B1(new_n258), .B2(new_n515), .ZN(new_n516));
  MUX2_X1   g0316(.A(G257), .B(G264), .S(G1698), .Z(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n258), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(G270), .B1(new_n474), .B2(new_n475), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n478), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n514), .A2(KEYINPUT21), .A3(G169), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n505), .B1(new_n506), .B2(new_n504), .ZN(new_n524));
  INV_X1    g0324(.A(new_n513), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n511), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n522), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n520), .A2(new_n295), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n514), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n520), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n526), .B1(new_n531), .B2(new_n343), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n532), .A2(KEYINPUT82), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n532), .A2(KEYINPUT82), .B1(G190), .B2(new_n531), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n215), .B1(new_n323), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n224), .A3(new_n442), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n255), .A2(new_n257), .A3(new_n215), .A4(G68), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n288), .B2(new_n224), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n280), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n447), .A2(new_n361), .ZN(new_n545));
  INV_X1    g0345(.A(new_n361), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n503), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n231), .A2(new_n252), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n223), .A2(G1698), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n251), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n254), .A2(new_n504), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n266), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n475), .A2(G250), .ZN(new_n555));
  INV_X1    g0355(.A(new_n477), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n277), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n477), .B1(new_n475), .B2(G250), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n549), .A2(new_n550), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n552), .B1(new_n560), .B2(new_n251), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n295), .B(new_n559), .C1(new_n561), .C2(new_n266), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n548), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G200), .B1(new_n554), .B2(new_n557), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n447), .A2(G87), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n543), .A2(new_n280), .B1(new_n503), .B2(new_n546), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G190), .B(new_n559), .C1(new_n561), .C2(new_n266), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n565), .A2(new_n568), .A3(new_n567), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT81), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G264), .B1(new_n474), .B2(new_n475), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n225), .B2(G1698), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n251), .B1(G33), .B2(G294), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n478), .C1(new_n266), .C2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n405), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G200), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n215), .A2(G107), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT85), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n442), .A2(G20), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT23), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n582), .C2(new_n583), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(new_n215), .B2(new_n552), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n255), .A2(new_n257), .A3(new_n215), .A4(G87), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n591), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n594), .A3(KEYINPUT24), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n280), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT25), .B1(new_n283), .B2(G107), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n283), .A2(KEYINPUT25), .A3(G107), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n506), .C2(new_n442), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n581), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n579), .A2(new_n277), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(G179), .B2(new_n579), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n599), .B2(new_n603), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n535), .A2(new_n574), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n437), .A2(new_n502), .A3(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n428), .A2(new_n423), .ZN(new_n611));
  INV_X1    g0411(.A(new_n342), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n349), .B2(new_n374), .ZN(new_n613));
  INV_X1    g0413(.A(new_n415), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n303), .A2(new_n305), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n297), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n565), .A2(new_n568), .A3(new_n570), .A4(new_n567), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n563), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n604), .B(new_n620), .C1(new_n607), .C2(new_n530), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n502), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n479), .B1(new_n489), .B2(new_n496), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n481), .B1(G200), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g0424(.A(G179), .B(new_n483), .C1(new_n484), .C2(new_n486), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n444), .A2(new_n448), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n483), .B1(new_n267), .B2(new_n495), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(G169), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT80), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n621), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(KEYINPUT87), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n497), .A2(new_n499), .A3(new_n620), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n635), .A3(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n630), .A4(new_n574), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n563), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n617), .B1(new_n437), .B2(new_n645), .ZN(G369));
  AND2_X1   g0446(.A1(new_n599), .A2(new_n603), .ZN(new_n647));
  XOR2_X1   g0447(.A(KEYINPUT89), .B(KEYINPUT27), .Z(new_n648));
  NOR3_X1   g0448(.A1(new_n208), .A2(G1), .A3(G20), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n604), .B1(new_n647), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n608), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n607), .A2(new_n654), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n530), .A2(new_n654), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n654), .A2(new_n526), .ZN(new_n663));
  MUX2_X1   g0463(.A(new_n535), .B(new_n530), .S(new_n663), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n656), .A2(new_n661), .B1(new_n607), .B2(new_n654), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(G399));
  NOR2_X1   g0469(.A1(new_n539), .A2(G116), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT90), .Z(new_n671));
  NOR2_X1   g0471(.A1(new_n211), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n220), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(new_n654), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n622), .A2(new_n633), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n636), .A2(new_n635), .A3(new_n637), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n638), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n564), .B1(new_n681), .B2(new_n642), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n629), .A2(new_n637), .A3(new_n630), .A4(new_n574), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n564), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT93), .B1(new_n502), .B2(new_n621), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n631), .A2(new_n690), .A3(new_n632), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n654), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n685), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n559), .B1(new_n561), .B2(new_n266), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n520), .A2(new_n295), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n579), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT92), .B1(new_n487), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n623), .A2(new_n701), .A3(new_n579), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n575), .B1(new_n578), .B2(new_n266), .ZN(new_n704));
  NOR4_X1   g0504(.A1(new_n520), .A2(new_n704), .A3(new_n697), .A4(new_n295), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n627), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n627), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n696), .B(new_n678), .C1(new_n703), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n609), .A2(new_n502), .A3(new_n678), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n678), .B1(new_n703), .B2(new_n710), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n695), .B1(G330), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n677), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n664), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n208), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n269), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n672), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n721), .A2(new_n665), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n210), .A2(G355), .A3(new_n251), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G116), .B2(new_n210), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n211), .A2(new_n251), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n220), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n246), .A2(new_n733), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n214), .B1(G20), .B2(new_n277), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n725), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n405), .A2(G20), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n343), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G283), .A2(new_n749), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n295), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n753), .B(new_n258), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n745), .A2(new_n295), .A3(new_n343), .ZN(new_n758));
  INV_X1    g0558(.A(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n215), .A2(new_n405), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n747), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n755), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n762), .B1(new_n515), .B2(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n215), .B1(new_n750), .B2(G190), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(G20), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT99), .B(G326), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n773), .A2(G294), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n768), .B1(new_n781), .B2(KEYINPUT100), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(KEYINPUT100), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n756), .A2(new_n202), .B1(new_n766), .B2(new_n228), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n778), .B2(G50), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT97), .B(G159), .Z(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n751), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n773), .A2(G97), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n258), .B1(new_n749), .B2(G107), .ZN(new_n792));
  INV_X1    g0592(.A(new_n764), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G87), .B1(new_n758), .B2(G68), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n782), .A2(new_n783), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n744), .B1(new_n796), .B2(new_n741), .ZN(new_n797));
  INV_X1    g0597(.A(new_n740), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n664), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n728), .A2(new_n799), .ZN(G396));
  NAND4_X1  g0600(.A1(new_n368), .A2(new_n373), .A3(new_n365), .A4(new_n654), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n357), .A2(new_n366), .B1(new_n365), .B2(new_n678), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n374), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n683), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n716), .A2(G330), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n725), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n741), .A2(new_n738), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n725), .B1(G77), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n804), .A2(new_n739), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n756), .A2(new_n504), .B1(new_n764), .B2(new_n442), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n251), .B(new_n814), .C1(G87), .C2(new_n749), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n778), .A2(G303), .ZN(new_n816));
  INV_X1    g0616(.A(new_n758), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n817), .A2(new_n818), .B1(new_n751), .B2(new_n754), .ZN(new_n819));
  INV_X1    g0619(.A(new_n766), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G294), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n816), .A3(new_n791), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n756), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(new_n787), .B1(new_n820), .B2(G143), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n284), .B2(new_n817), .C1(new_n777), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n749), .A2(G68), .B1(new_n793), .B2(G50), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n258), .B1(new_n752), .B2(G132), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n772), .C2(new_n228), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(KEYINPUT101), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n822), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n812), .B(new_n813), .C1(new_n741), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n809), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  XOR2_X1   g0637(.A(new_n440), .B(KEYINPUT102), .Z(new_n838));
  INV_X1    g0638(.A(KEYINPUT35), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n504), .B(new_n217), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT36), .Z(new_n842));
  OR3_X1    g0642(.A1(new_n220), .A2(new_n202), .A3(new_n382), .ZN(new_n843));
  INV_X1    g0643(.A(G50), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n269), .B(G13), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n430), .A2(new_n416), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n416), .A2(new_n653), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n411), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n416), .A2(KEYINPUT104), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n391), .A2(new_n856), .A3(new_n393), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n430), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n653), .A3(new_n857), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n411), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n854), .B1(KEYINPUT37), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n859), .B1(new_n415), .B2(new_n432), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n859), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n433), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n853), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n347), .B2(new_n654), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n320), .A2(KEYINPUT103), .A3(new_n678), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n342), .A2(new_n349), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n320), .B(new_n678), .C1(new_n334), .C2(new_n341), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n803), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n609), .A2(new_n502), .A3(new_n678), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n876), .B(new_n711), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n848), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n411), .A2(new_n850), .A3(new_n852), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n851), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n852), .B1(new_n415), .B2(new_n611), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n849), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n868), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n885), .A2(new_n716), .A3(KEYINPUT40), .A4(new_n876), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n880), .A2(new_n436), .A3(new_n716), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n879), .B1(new_n868), .B2(new_n863), .ZN(new_n888));
  OAI211_X1 g0688(.A(G330), .B(new_n886), .C1(new_n888), .C2(KEYINPUT40), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n437), .A2(new_n806), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n695), .A2(new_n436), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n617), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n892), .B(new_n894), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n874), .A2(new_n875), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n654), .B(new_n804), .C1(new_n634), .C2(new_n644), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n801), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n869), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n428), .A2(new_n423), .A3(new_n652), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n342), .A2(new_n678), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n884), .A2(new_n868), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n863), .B2(new_n868), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n895), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n269), .B2(new_n722), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n895), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n847), .B1(new_n910), .B2(new_n911), .ZN(G367));
  NAND2_X1  g0712(.A1(new_n678), .A2(new_n626), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n625), .A2(new_n628), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n631), .A2(new_n913), .B1(new_n914), .B2(new_n678), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n667), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n608), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n500), .A2(new_n501), .ZN(new_n919));
  OR3_X1    g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n654), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n659), .A2(new_n661), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n923), .A2(KEYINPUT42), .A3(new_n502), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT42), .B1(new_n923), .B2(new_n502), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n921), .A2(new_n654), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n926), .B1(new_n929), .B2(new_n920), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT43), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT43), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n928), .B2(KEYINPUT106), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n928), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n568), .A2(new_n567), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n678), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n620), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n563), .B2(new_n937), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n928), .A2(KEYINPUT106), .A3(new_n933), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(KEYINPUT107), .B(new_n916), .C1(new_n940), .C2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT107), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n935), .B2(new_n939), .ZN(new_n946));
  INV_X1    g0746(.A(new_n916), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n914), .A2(new_n678), .ZN(new_n949));
  INV_X1    g0749(.A(new_n913), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n502), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n668), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n668), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n666), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n662), .A2(new_n665), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n667), .A2(new_n923), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n717), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n672), .B(KEYINPUT41), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n724), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n946), .B2(new_n947), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n944), .A2(new_n948), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n741), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n756), .A2(new_n844), .B1(new_n766), .B2(new_n284), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n258), .B(new_n967), .C1(G58), .C2(new_n793), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n778), .A2(G143), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n773), .A2(G68), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n748), .A2(new_n202), .B1(new_n751), .B2(new_n825), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n787), .B2(new_n758), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G294), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n793), .A2(G116), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT46), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n258), .B1(new_n817), .B2(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n778), .A2(G311), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G97), .A2(new_n749), .B1(new_n752), .B2(G317), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n823), .A2(G283), .B1(new_n820), .B2(G303), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n772), .A2(new_n442), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n973), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n966), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n732), .A2(new_n242), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n743), .B1(new_n211), .B2(new_n361), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n726), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n798), .C2(new_n939), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n965), .A2(new_n991), .ZN(G387));
  INV_X1    g0792(.A(new_n960), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n658), .A2(new_n740), .ZN(new_n994));
  INV_X1    g0794(.A(new_n291), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT50), .B1(new_n995), .B2(G50), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n733), .C1(new_n230), .C2(new_n202), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n995), .A2(KEYINPUT50), .A3(G50), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n258), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n671), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n239), .A2(G45), .A3(new_n258), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n211), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n742), .B1(new_n442), .B2(new_n210), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n725), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n817), .A2(new_n995), .B1(new_n756), .B2(new_n230), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n258), .B(new_n1005), .C1(G97), .C2(new_n749), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n778), .A2(G159), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n773), .A2(new_n361), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n793), .A2(G77), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n284), .B2(new_n751), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G50), .B2(new_n820), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n823), .A2(G303), .B1(G311), .B2(new_n758), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n759), .B2(new_n766), .C1(new_n777), .C2(new_n765), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n773), .A2(G283), .B1(G294), .B2(new_n793), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT109), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT49), .Z(new_n1021));
  INV_X1    g0821(.A(new_n779), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n258), .B1(new_n748), .B2(new_n504), .C1(new_n751), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1012), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1004), .B1(new_n1024), .B2(new_n741), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n993), .A2(new_n724), .B1(new_n994), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n993), .A2(new_n806), .A3(new_n694), .A4(new_n685), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n672), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n717), .A2(new_n993), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(G393));
  XNOR2_X1  g0830(.A(new_n957), .B(new_n667), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n915), .A2(new_n740), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n742), .B1(new_n224), .B2(new_n210), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n249), .B2(new_n731), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n726), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT110), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n823), .A2(G294), .B1(G303), .B2(new_n758), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n818), .B2(new_n764), .C1(new_n765), .C2(new_n751), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n251), .B(new_n1038), .C1(G107), .C2(new_n749), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n777), .A2(new_n759), .B1(new_n754), .B2(new_n766), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT52), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n504), .C2(new_n772), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  INV_X1    g0844(.A(G159), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n777), .A2(new_n284), .B1(new_n1045), .B2(new_n766), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT51), .Z(new_n1047));
  NOR2_X1   g0847(.A1(new_n764), .A2(new_n230), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n251), .B1(new_n748), .B2(new_n538), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G143), .C2(new_n752), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n817), .A2(new_n844), .B1(new_n995), .B2(new_n756), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n773), .A2(G77), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1043), .A2(new_n1044), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1036), .B1(new_n1056), .B2(new_n741), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1031), .A2(new_n724), .B1(new_n1032), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1031), .B1(new_n717), .B2(new_n993), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n672), .B1(new_n1027), .B2(new_n958), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(G390));
  NAND4_X1  g0861(.A1(new_n716), .A2(G330), .A3(new_n804), .A4(new_n896), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(KEYINPUT114), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n802), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n375), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n692), .A2(new_n654), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n801), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT112), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(KEYINPUT112), .A3(new_n801), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n896), .B(KEYINPUT113), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n902), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n801), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n683), .B2(new_n804), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1076), .B2(new_n897), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n904), .A2(new_n905), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1073), .A2(new_n885), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1062), .A2(KEYINPUT114), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n906), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1063), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1078), .B1(new_n899), .B2(new_n902), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1066), .A2(KEYINPUT112), .A3(new_n801), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT112), .B1(new_n1066), .B2(new_n801), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n1071), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n885), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1063), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1081), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n724), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1078), .A2(new_n738), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n726), .B1(new_n995), .B2(new_n810), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n773), .A2(G159), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  AOI21_X1  g0897(.A(new_n258), .B1(new_n823), .B2(new_n1097), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n284), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT53), .B1(new_n764), .B2(new_n284), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n820), .A2(G132), .B1(new_n758), .B2(G137), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1102), .B1(new_n844), .B2(new_n748), .C1(new_n1103), .C2(new_n751), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(G128), .C2(new_n778), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n823), .A2(G97), .B1(G107), .B2(new_n758), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n504), .B2(new_n766), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n251), .B1(new_n793), .B2(G87), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n230), .B2(new_n748), .C1(new_n974), .C2(new_n751), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(G283), .C2(new_n778), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1096), .A2(new_n1105), .B1(new_n1110), .B2(new_n1053), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1094), .B(new_n1095), .C1(new_n966), .C2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n894), .A2(new_n891), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n716), .A2(G330), .A3(new_n804), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n897), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1062), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1076), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1071), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n1062), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1082), .A2(new_n1122), .A3(new_n1091), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n672), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1093), .B(new_n1112), .C1(new_n1124), .C2(new_n1125), .ZN(G378));
  NOR2_X1   g0926(.A1(G33), .A2(G41), .ZN(new_n1127));
  INV_X1    g0927(.A(G124), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1127), .B1(new_n751), .B2(new_n1128), .C1(new_n788), .C2(new_n748), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G128), .A2(new_n820), .B1(new_n793), .B2(new_n1097), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n823), .A2(G137), .B1(G132), .B2(new_n758), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n284), .B2(new_n772), .C1(new_n777), .C2(new_n1103), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1133), .B2(KEYINPUT59), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(KEYINPUT59), .B2(new_n1133), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT58), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n251), .A2(G41), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n817), .B2(new_n224), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n752), .A2(G283), .B1(new_n820), .B2(G107), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n749), .A2(G58), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1009), .A3(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1138), .B(new_n1141), .C1(new_n361), .C2(new_n823), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n970), .C1(new_n504), .C2(new_n777), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1137), .A2(G50), .A3(new_n1127), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT115), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1135), .B1(new_n1136), .B2(new_n1143), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n741), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1149), .B(new_n725), .C1(G50), .C2(new_n811), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n306), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n294), .A2(new_n653), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT116), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1155), .B2(new_n738), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT117), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n906), .A2(new_n901), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1076), .A2(new_n870), .A3(new_n897), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n889), .A2(new_n1155), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1151), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n306), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n306), .A2(new_n1163), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1164), .A2(new_n1154), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1154), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(new_n880), .A3(G330), .A4(new_n886), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1161), .B(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1157), .B1(new_n1171), .B2(new_n724), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n893), .B(new_n617), .C1(new_n437), .C2(new_n806), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1120), .B2(new_n1118), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1079), .A2(new_n1063), .A3(new_n1081), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1089), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1113), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1171), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1092), .B2(new_n1121), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1170), .A2(new_n907), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n908), .A2(new_n1169), .A3(new_n1162), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT57), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n672), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1172), .B1(new_n1179), .B2(new_n1185), .ZN(G375));
  NAND3_X1  g0986(.A1(new_n1173), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1122), .A2(new_n962), .A3(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n817), .A2(new_n504), .B1(new_n751), .B2(new_n515), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n251), .B(new_n1189), .C1(G77), .C2(new_n749), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n778), .A2(G294), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n756), .A2(new_n442), .B1(new_n764), .B2(new_n224), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G283), .B2(new_n820), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1008), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n823), .A2(G150), .B1(new_n820), .B2(G137), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1195), .A2(new_n251), .A3(new_n1140), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n758), .A2(new_n1097), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1045), .B2(new_n764), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G128), .B2(new_n752), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n773), .A2(G50), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n778), .A2(G132), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1196), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1194), .A2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n725), .B1(G68), .B2(new_n811), .C1(new_n1203), .C2(new_n966), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1071), .B2(new_n738), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n723), .B(KEYINPUT119), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1121), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1188), .A2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(KEYINPUT121), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G375), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G378), .ZN(new_n1211));
  OAI211_X1 g1011(.A(KEYINPUT57), .B(new_n1183), .C1(new_n1125), .C2(new_n1173), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1170), .B(new_n1160), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1177), .B2(new_n1113), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1212), .B(new_n672), .C1(new_n1214), .C2(KEYINPUT57), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1210), .A2(new_n1211), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G387), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G381), .A2(G390), .ZN(new_n1220));
  INV_X1    g1020(.A(G396), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n1026), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G384), .A2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1224), .ZN(G407));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G343), .C2(new_n1217), .ZN(G409));
  NAND2_X1  g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1222), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(G390), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1229), .A2(new_n965), .A3(new_n991), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n965), .B2(new_n991), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT123), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1172), .C1(new_n1179), .C2(new_n1185), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1206), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1157), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT122), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1171), .B(new_n962), .C1(new_n1125), .C2(new_n1173), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT122), .B1(new_n1239), .B2(new_n1157), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1211), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1237), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1187), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1187), .A2(new_n1252), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n672), .A3(new_n1122), .A4(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1207), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(G384), .B1(new_n1255), .B2(new_n1207), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1248), .A2(new_n1251), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(KEYINPUT61), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(KEYINPUT61), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1236), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G2897), .B(new_n1250), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1258), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1250), .A2(G2897), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1256), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1248), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1250), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1274), .B(new_n1277), .C1(new_n1275), .C2(new_n1250), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1260), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1251), .A4(new_n1259), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1269), .A2(new_n1276), .B1(new_n1235), .B2(new_n1283), .ZN(G405));
  AND3_X1   g1084(.A1(new_n1271), .A2(KEYINPUT125), .A3(new_n1256), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1237), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1215), .B2(new_n1172), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1211), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1271), .A2(KEYINPUT125), .A3(new_n1256), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1237), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1289), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT127), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1288), .A2(new_n1292), .A3(new_n1289), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1234), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1294), .A2(new_n1299), .A3(new_n1234), .A4(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(G402));
endmodule


