//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n188), .B(G146), .C1(KEYINPUT16), .C2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n198), .B(KEYINPUT74), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT75), .B1(new_n194), .B2(G128), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n195), .A3(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT76), .B(G110), .Z(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n191), .B(new_n193), .C1(new_n201), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n199), .A2(new_n200), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G110), .ZN(new_n210));
  INV_X1    g024(.A(new_n191), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n187), .B2(KEYINPUT16), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n218), .B(KEYINPUT77), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n216), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT69), .B(G902), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(KEYINPUT78), .B2(KEYINPUT25), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  OAI21_X1  g043(.A(G217), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT73), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n228), .B(new_n232), .C1(new_n226), .C2(new_n224), .ZN(new_n233));
  INV_X1    g047(.A(new_n222), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n232), .A2(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n239), .B2(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n241), .A2(new_n242), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n243), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n247), .B2(new_n240), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n192), .A2(G143), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT64), .A3(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(G128), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(KEYINPUT1), .A3(new_n196), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n251), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G143), .B(G146), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n196), .B1(new_n253), .B2(new_n254), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n257), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n267), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n250), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G116), .B(G119), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT65), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT2), .B(G113), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n246), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT0), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n265), .B1(new_n281), .B2(new_n196), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT0), .B(G128), .Z(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n265), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n269), .A2(new_n277), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n261), .A2(new_n263), .A3(new_n251), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT66), .B1(new_n267), .B2(new_n262), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n249), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n285), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n276), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n291), .A3(KEYINPUT68), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n293), .B(new_n276), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n285), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n289), .B2(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n298), .A3(new_n277), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G237), .A2(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G210), .ZN(new_n303));
  INV_X1    g117(.A(G101), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n295), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n223), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT70), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n285), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n250), .B1(new_n267), .B2(new_n262), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n285), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n276), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n286), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n320), .B2(new_n307), .ZN(new_n321));
  INV_X1    g135(.A(new_n286), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n277), .B1(new_n285), .B2(new_n315), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT28), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n301), .A2(new_n324), .A3(new_n308), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n312), .A2(new_n313), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G472), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT71), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n286), .A3(new_n308), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n319), .A2(KEYINPUT31), .A3(new_n286), .A4(new_n308), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n301), .A2(new_n324), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n307), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G472), .A2(G902), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n337), .A2(KEYINPUT32), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT32), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n313), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n311), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n325), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G472), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n347), .A4(new_n341), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n238), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G214), .B1(G237), .B2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n355), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G104), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G101), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(G101), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n356), .A2(new_n359), .A3(new_n304), .A4(new_n360), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n276), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n355), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n358), .A2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n271), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n194), .A3(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G113), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n275), .B(new_n372), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G110), .B(G122), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n377), .A3(new_n379), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n284), .A2(KEYINPUT84), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT84), .B1(new_n284), .B2(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n261), .A2(new_n263), .A3(new_n384), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT85), .B(G224), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n388), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n378), .A2(new_n393), .A3(new_n380), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G902), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT7), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n388), .A2(new_n397), .A3(new_n391), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n388), .B1(new_n397), .B2(new_n391), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n379), .B(KEYINPUT8), .Z(new_n400));
  AND2_X1   g214(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n275), .B1(new_n401), .B2(new_n376), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n372), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n275), .B1(new_n374), .B2(new_n376), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n372), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n398), .A2(new_n399), .A3(new_n382), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n396), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n395), .A2(new_n396), .A3(new_n408), .A4(new_n406), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n354), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G469), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT10), .B(new_n372), .C1(new_n264), .C2(new_n268), .ZN(new_n417));
  INV_X1    g231(.A(new_n280), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n366), .A2(new_n284), .A3(new_n363), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT10), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n256), .A2(new_n259), .A3(G128), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT1), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n253), .A2(G128), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n260), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n424), .B2(new_n371), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n417), .A2(new_n426), .A3(KEYINPUT80), .A4(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n217), .A2(G227), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n432), .B(new_n433), .Z(new_n434));
  AOI21_X1  g248(.A(new_n416), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  AOI211_X1 g250(.A(KEYINPUT82), .B(new_n436), .C1(new_n429), .C2(new_n430), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n372), .A2(new_n267), .A3(new_n262), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n424), .A2(new_n371), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n280), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n418), .B2(KEYINPUT81), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n435), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n417), .A2(new_n426), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n429), .A2(new_n430), .B1(new_n280), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(new_n434), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n280), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n419), .A2(new_n425), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n371), .B1(new_n287), .B2(new_n288), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(KEYINPUT10), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT80), .B1(new_n452), .B2(new_n418), .ZN(new_n453));
  INV_X1    g267(.A(new_n430), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT83), .A3(new_n436), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n415), .B(new_n311), .C1(new_n444), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(G469), .A2(G902), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n453), .A2(new_n454), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n436), .B1(new_n460), .B2(new_n443), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n447), .A2(new_n434), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n458), .B(new_n459), .C1(new_n415), .C2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n465));
  AOI21_X1  g279(.A(G143), .B1(new_n302), .B2(G214), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT18), .B(G131), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n302), .A2(G214), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n252), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n384), .A2(G140), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n190), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n193), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n193), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n473), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(KEYINPUT19), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT19), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n190), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n482), .A2(new_n483), .A3(new_n192), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n191), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n465), .B2(new_n466), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n469), .A2(new_n470), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(G131), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n242), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n487), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n482), .A2(new_n485), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n483), .B1(new_n497), .B2(new_n192), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n481), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(G113), .B(G122), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT90), .B(G104), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT91), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n211), .A2(new_n214), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n493), .A2(new_n495), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(KEYINPUT17), .ZN(new_n509));
  INV_X1    g323(.A(new_n481), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n489), .A2(new_n492), .B1(new_n242), .B2(new_n494), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n513), .A2(new_n498), .A3(new_n487), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n503), .C1(new_n514), .C2(new_n481), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n505), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G475), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n396), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n520), .A3(new_n517), .A4(new_n396), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n511), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n396), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G475), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT9), .B(G234), .Z(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G217), .A3(new_n217), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT13), .B1(new_n252), .B2(G128), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n252), .A2(G128), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n252), .A2(KEYINPUT13), .A3(G128), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n196), .B2(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n196), .A2(G143), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G134), .ZN(new_n540));
  XOR2_X1   g354(.A(G116), .B(G122), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(G107), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n252), .A2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n537), .A3(new_n239), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT93), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n547));
  INV_X1    g361(.A(G116), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT14), .A3(G122), .ZN(new_n549));
  OAI211_X1 g363(.A(G107), .B(new_n549), .C1(new_n541), .C2(KEYINPUT14), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n537), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G134), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n550), .B(new_n553), .C1(G107), .C2(new_n541), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n546), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n547), .B1(new_n546), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n529), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n546), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n559));
  INV_X1    g373(.A(new_n529), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n546), .A2(new_n554), .A3(new_n547), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n311), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(KEYINPUT15), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n217), .A2(G952), .ZN(new_n572));
  NAND2_X1  g386(.A1(G234), .A2(G237), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT96), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT21), .B(G898), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n223), .A2(G953), .A3(new_n573), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n527), .A2(new_n571), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G221), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n528), .B2(new_n396), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n414), .A2(new_n464), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n352), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT97), .B(G101), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G3));
  NAND2_X1  g404(.A1(new_n337), .A2(new_n311), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n337), .A2(new_n338), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n464), .A3(new_n237), .A4(new_n585), .ZN(new_n596));
  INV_X1    g410(.A(new_n412), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT33), .B1(new_n557), .B2(new_n562), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n602), .A2(KEYINPUT98), .A3(G478), .A4(new_n311), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n563), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(G478), .A3(new_n311), .A4(new_n599), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n564), .A2(new_n567), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n527), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n581), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n527), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n581), .B(KEYINPUT99), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n571), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT100), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n598), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  NOR2_X1   g439(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n216), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n235), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT103), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n233), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n592), .A2(new_n630), .A3(new_n593), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n592), .A2(new_n630), .A3(KEYINPUT104), .A4(new_n593), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n586), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT37), .B(G110), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  NAND2_X1  g452(.A1(new_n350), .A2(new_n351), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n464), .A2(new_n585), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n616), .A2(new_n571), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n576), .B1(new_n580), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n630), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n597), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n639), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n644), .B(KEYINPUT39), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n640), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n527), .A2(new_n571), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n330), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n292), .A2(new_n307), .A3(new_n294), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(KEYINPUT105), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(KEYINPUT105), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n396), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n341), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n410), .A2(new_n411), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT38), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n353), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n656), .A2(new_n630), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT106), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(new_n644), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n527), .A2(new_n610), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n639), .A2(new_n641), .A3(new_n647), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  OAI21_X1  g488(.A(new_n311), .B1(new_n444), .B2(new_n457), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(KEYINPUT107), .A3(new_n458), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n678), .A3(G469), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n597), .B(new_n584), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n639), .A2(new_n237), .A3(new_n612), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n639), .A2(new_n620), .A3(new_n237), .A4(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT108), .B(G116), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G18));
  NAND4_X1  g500(.A1(new_n639), .A2(new_n582), .A3(new_n630), .A4(new_n680), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(G119), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G21));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n295), .A2(new_n690), .A3(new_n301), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n307), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n690), .B1(new_n295), .B2(new_n301), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n334), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n338), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n237), .A2(new_n592), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT111), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n680), .A2(new_n697), .A3(new_n618), .A4(new_n655), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  XNOR2_X1  g513(.A(new_n671), .B(KEYINPUT112), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n592), .A2(new_n695), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n680), .A3(new_n630), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n461), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT113), .B(new_n436), .C1(new_n460), .C2(new_n443), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(G469), .A3(new_n462), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n458), .A2(new_n459), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n664), .A2(new_n354), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n585), .A3(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n639), .A3(new_n237), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n671), .B(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n711), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n348), .A2(new_n237), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT42), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n242), .ZN(G33));
  NAND4_X1  g535(.A1(new_n639), .A2(new_n237), .A3(new_n645), .A4(new_n716), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  NAND4_X1  g537(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n462), .A4(new_n707), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n463), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(G469), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n459), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n458), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT46), .B1(new_n727), .B2(new_n459), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n585), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n731), .A2(new_n651), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n710), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n616), .A2(new_n610), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n594), .A3(new_n630), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n733), .B(new_n740), .C1(new_n739), .C2(new_n738), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  OR2_X1    g556(.A1(new_n731), .A2(KEYINPUT114), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n731), .A2(KEYINPUT114), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n748), .A3(new_n744), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n639), .A2(new_n671), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n238), .A3(new_n710), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G140), .ZN(G42));
  NAND2_X1  g567(.A1(new_n677), .A2(new_n679), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT49), .Z(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n663), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n665), .A2(new_n735), .A3(new_n584), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n237), .A3(new_n353), .A4(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n737), .A2(new_n576), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n697), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n585), .B1(new_n677), .B2(new_n679), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n710), .B(new_n761), .C1(new_n750), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n754), .A2(new_n585), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n665), .A2(new_n353), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n765), .A2(KEYINPUT50), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n764), .A2(new_n734), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n759), .A2(new_n772), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n773), .A2(new_n646), .A3(new_n701), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n763), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n763), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n663), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n772), .A2(new_n237), .A3(new_n576), .A4(new_n778), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n779), .A2(new_n527), .A3(new_n610), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n763), .A2(new_n771), .A3(new_n780), .A4(new_n774), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n781), .A2(new_n784), .A3(new_n572), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n761), .A2(new_n680), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n681), .A2(new_n687), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n684), .A2(new_n698), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n642), .A2(new_n611), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n414), .A3(new_n618), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n596), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n792), .B(new_n636), .C1(new_n352), .C2(new_n587), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n722), .A2(new_n713), .A3(new_n719), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n527), .A2(new_n571), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n670), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n640), .B(new_n797), .C1(new_n350), .C2(new_n351), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n709), .A2(new_n585), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n700), .A2(new_n701), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n630), .B(new_n710), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n799), .A2(new_n630), .A3(new_n644), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n655), .A2(new_n412), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n663), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n673), .A2(new_n649), .A3(new_n703), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n640), .B1(new_n350), .B2(new_n351), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n412), .A2(new_n754), .A3(new_n585), .A4(new_n630), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n809), .A2(new_n648), .B1(new_n810), .B2(new_n702), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n673), .A4(new_n806), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n681), .A2(new_n684), .A3(new_n687), .A4(new_n698), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n793), .A3(new_n795), .A4(new_n801), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n808), .A2(new_n813), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n787), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n681), .A2(new_n684), .A3(new_n687), .A4(new_n698), .ZN(new_n826));
  INV_X1    g640(.A(new_n636), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n588), .B(new_n827), .C1(new_n596), .C2(new_n791), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n795), .A2(new_n801), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n823), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n785), .A2(new_n786), .A3(new_n825), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n779), .A2(new_n611), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n773), .A2(new_n718), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT48), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(G952), .A2(G953), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n758), .B1(new_n838), .B2(new_n839), .ZN(G75));
  NAND2_X1  g654(.A1(new_n383), .A2(new_n394), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n392), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT55), .Z(new_n843));
  AOI21_X1  g657(.A(KEYINPUT116), .B1(new_n831), .B2(new_n823), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n830), .A2(new_n829), .A3(new_n808), .A4(new_n813), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n787), .B1(new_n845), .B2(new_n819), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n223), .B(new_n409), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n843), .B1(new_n848), .B2(KEYINPUT56), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n217), .A2(G952), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  INV_X1    g666(.A(new_n843), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n849), .A2(KEYINPUT118), .A3(new_n851), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(G51));
  INV_X1    g673(.A(new_n727), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n223), .B(new_n860), .C1(new_n844), .C2(new_n846), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n459), .B(KEYINPUT57), .Z(new_n863));
  AOI21_X1  g677(.A(new_n822), .B1(new_n821), .B2(new_n824), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n844), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n444), .A2(new_n457), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT119), .B1(new_n868), .B2(new_n850), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  INV_X1    g684(.A(new_n867), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n844), .B2(new_n846), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n825), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(new_n863), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n870), .B(new_n851), .C1(new_n874), .C2(new_n862), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n875), .ZN(G54));
  AOI21_X1  g690(.A(new_n311), .B1(new_n821), .B2(new_n824), .ZN(new_n877));
  AND2_X1   g691(.A1(KEYINPUT58), .A2(G475), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(KEYINPUT120), .A3(new_n516), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n223), .B(new_n878), .C1(new_n844), .C2(new_n846), .ZN(new_n881));
  INV_X1    g695(.A(new_n516), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n850), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(G60));
  AND2_X1   g704(.A1(new_n825), .A2(new_n833), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT59), .Z(new_n893));
  OAI22_X1  g707(.A1(new_n891), .A2(new_n893), .B1(new_n600), .B2(new_n601), .ZN(new_n894));
  INV_X1    g708(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n873), .A2(new_n602), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n851), .A3(new_n896), .ZN(G63));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT60), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n821), .B2(new_n824), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n850), .B1(new_n900), .B2(new_n627), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n234), .B2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(G66));
  OAI21_X1  g718(.A(G953), .B1(new_n578), .B2(new_n390), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n794), .B(KEYINPUT122), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n841), .B1(G898), .B2(new_n217), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(G69));
  NAND2_X1  g723(.A1(new_n314), .A2(new_n318), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n497), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n652), .A2(new_n734), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n352), .A3(new_n790), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n752), .A2(new_n741), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT106), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n667), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n811), .A2(new_n673), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n918), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n668), .A2(KEYINPUT62), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n914), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n922), .B2(G953), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n733), .A2(new_n237), .A3(new_n348), .A4(new_n805), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n752), .A2(new_n741), .A3(new_n920), .A4(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n795), .B(KEYINPUT125), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n911), .B1(new_n929), .B2(new_n217), .ZN(new_n930));
  NAND2_X1  g744(.A1(G900), .A2(G953), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT124), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT123), .B(new_n911), .C1(new_n922), .C2(G953), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n925), .A2(new_n937), .A3(new_n932), .A4(new_n933), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G72));
  NAND2_X1  g753(.A1(new_n320), .A2(new_n307), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n330), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n307), .B1(new_n927), .B2(new_n928), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n906), .B(new_n942), .C1(new_n922), .C2(new_n307), .ZN(new_n943));
  XOR2_X1   g757(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n328), .A2(new_n396), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT127), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n941), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n832), .A2(new_n941), .A3(new_n946), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n850), .A3(new_n949), .ZN(G57));
endmodule


