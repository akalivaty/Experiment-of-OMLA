

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  INV_X1 U325 ( .A(KEYINPUT94), .ZN(n365) );
  XNOR2_X1 U326 ( .A(n366), .B(n365), .ZN(n370) );
  XNOR2_X1 U327 ( .A(n327), .B(n326), .ZN(n328) );
  NOR2_X1 U328 ( .A1(n504), .A2(n518), .ZN(n455) );
  XOR2_X1 U329 ( .A(KEYINPUT70), .B(n442), .Z(n293) );
  XOR2_X1 U330 ( .A(n398), .B(n452), .Z(n294) );
  XOR2_X1 U331 ( .A(n447), .B(n446), .Z(n295) );
  XOR2_X1 U332 ( .A(KEYINPUT45), .B(n465), .Z(n296) );
  INV_X1 U333 ( .A(KEYINPUT91), .ZN(n324) );
  XNOR2_X1 U334 ( .A(n325), .B(n324), .ZN(n326) );
  INV_X1 U335 ( .A(n585), .ZN(n422) );
  INV_X1 U336 ( .A(KEYINPUT11), .ZN(n392) );
  OR2_X1 U337 ( .A1(n589), .A2(n422), .ZN(n423) );
  XNOR2_X1 U338 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U339 ( .A(n448), .B(n295), .ZN(n449) );
  XNOR2_X1 U340 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U341 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U342 ( .A1(n532), .A2(n474), .ZN(n573) );
  NOR2_X1 U343 ( .A1(n484), .A2(n526), .ZN(n545) );
  XOR2_X1 U344 ( .A(n399), .B(n398), .Z(n556) );
  XNOR2_X1 U345 ( .A(n349), .B(n348), .ZN(n536) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n478) );
  XNOR2_X1 U347 ( .A(n485), .B(G120GAT), .ZN(n486) );
  XNOR2_X1 U348 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n298) );
  XNOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n299), .B(G85GAT), .Z(n301) );
  XOR2_X1 U353 ( .A(G1GAT), .B(G127GAT), .Z(n407) );
  XNOR2_X1 U354 ( .A(G148GAT), .B(n407), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G134GAT), .Z(n397) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n302), .B(G120GAT), .ZN(n341) );
  XOR2_X1 U359 ( .A(n397), .B(n341), .Z(n304) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U362 ( .A(n306), .B(n305), .Z(n317) );
  XOR2_X1 U363 ( .A(G155GAT), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(KEYINPUT84), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U366 ( .A(KEYINPUT83), .B(KEYINPUT2), .Z(n310) );
  XNOR2_X1 U367 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n354) );
  XOR2_X1 U370 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n314) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n354), .B(n315), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n372) );
  XNOR2_X1 U375 ( .A(KEYINPUT27), .B(KEYINPUT93), .ZN(n332) );
  XOR2_X1 U376 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n319) );
  XNOR2_X1 U377 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(G169GAT), .B(n320), .Z(n345) );
  XOR2_X1 U380 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G92GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n321), .B(G64GAT), .ZN(n452) );
  NAND2_X1 U383 ( .A1(G226GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n294), .B(n322), .ZN(n327) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n323), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U387 ( .A(n355), .B(KEYINPUT92), .ZN(n325) );
  XOR2_X1 U388 ( .A(G8GAT), .B(G183GAT), .Z(n405) );
  XOR2_X1 U389 ( .A(n328), .B(n405), .Z(n330) );
  XNOR2_X1 U390 ( .A(G204GAT), .B(G218GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U392 ( .A(n345), .B(n331), .Z(n471) );
  XOR2_X1 U393 ( .A(n332), .B(n471), .Z(n373) );
  XOR2_X1 U394 ( .A(G183GAT), .B(KEYINPUT80), .Z(n334) );
  XNOR2_X1 U395 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n349) );
  XOR2_X1 U397 ( .A(G134GAT), .B(G190GAT), .Z(n336) );
  XNOR2_X1 U398 ( .A(G43GAT), .B(G99GAT), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U400 ( .A(KEYINPUT20), .B(G71GAT), .Z(n338) );
  XNOR2_X1 U401 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U403 ( .A(n340), .B(n339), .Z(n347) );
  XOR2_X1 U404 ( .A(n341), .B(G176GAT), .Z(n343) );
  NAND2_X1 U405 ( .A1(G227GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U409 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n352) );
  INV_X1 U410 ( .A(G106GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n363) );
  XOR2_X1 U414 ( .A(G50GAT), .B(G218GAT), .Z(n391) );
  XOR2_X1 U415 ( .A(n355), .B(n391), .Z(n357) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n358), .B(KEYINPUT24), .Z(n361) );
  XNOR2_X1 U419 ( .A(G78GAT), .B(G204GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(G148GAT), .ZN(n445) );
  XNOR2_X1 U421 ( .A(n445), .B(KEYINPUT23), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n475) );
  NOR2_X1 U424 ( .A1(n536), .A2(n475), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n364), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U426 ( .A1(n373), .A2(n572), .ZN(n366) );
  NAND2_X1 U427 ( .A1(n471), .A2(n536), .ZN(n367) );
  NAND2_X1 U428 ( .A1(n475), .A2(n367), .ZN(n368) );
  XNOR2_X1 U429 ( .A(KEYINPUT25), .B(n368), .ZN(n369) );
  NOR2_X1 U430 ( .A1(n370), .A2(n369), .ZN(n371) );
  NOR2_X1 U431 ( .A1(n372), .A2(n371), .ZN(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT90), .B(n372), .ZN(n532) );
  NAND2_X1 U433 ( .A1(n532), .A2(n373), .ZN(n481) );
  XNOR2_X1 U434 ( .A(n475), .B(KEYINPUT66), .ZN(n374) );
  XOR2_X1 U435 ( .A(n374), .B(KEYINPUT28), .Z(n526) );
  OR2_X1 U436 ( .A1(n526), .A2(n536), .ZN(n375) );
  NOR2_X1 U437 ( .A1(n481), .A2(n375), .ZN(n376) );
  NOR2_X1 U438 ( .A1(n377), .A2(n376), .ZN(n490) );
  INV_X1 U439 ( .A(KEYINPUT36), .ZN(n400) );
  XOR2_X1 U440 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n379) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n386) );
  INV_X1 U443 ( .A(KEYINPUT71), .ZN(n380) );
  NAND2_X1 U444 ( .A1(n380), .A2(G85GAT), .ZN(n383) );
  INV_X1 U445 ( .A(G85GAT), .ZN(n381) );
  NAND2_X1 U446 ( .A1(n381), .A2(KEYINPUT71), .ZN(n382) );
  NAND2_X1 U447 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(G106GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n442) );
  XOR2_X1 U450 ( .A(n386), .B(n442), .Z(n390) );
  XOR2_X1 U451 ( .A(G43GAT), .B(KEYINPUT7), .Z(n388) );
  XNOR2_X1 U452 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n439) );
  XNOR2_X1 U454 ( .A(n439), .B(G162GAT), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n391), .B(G92GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n556), .ZN(n589) );
  XNOR2_X1 U459 ( .A(G22GAT), .B(G15GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n401), .B(KEYINPUT69), .ZN(n426) );
  XOR2_X1 U461 ( .A(n426), .B(KEYINPUT75), .Z(n403) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U464 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U465 ( .A(G71GAT), .B(G57GAT), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT13), .ZN(n444) );
  XNOR2_X1 U467 ( .A(n407), .B(n444), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U469 ( .A(G64GAT), .B(G211GAT), .Z(n411) );
  XNOR2_X1 U470 ( .A(G155GAT), .B(G78GAT), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U472 ( .A(n413), .B(n412), .Z(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT76), .B(KEYINPUT73), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT78), .B(KEYINPUT74), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n585) );
  OR2_X1 U481 ( .A1(n490), .A2(n423), .ZN(n425) );
  XOR2_X1 U482 ( .A(KEYINPUT37), .B(KEYINPUT98), .Z(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n504) );
  XOR2_X1 U484 ( .A(G29GAT), .B(n426), .Z(n428) );
  NAND2_X1 U485 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n429), .B(G36GAT), .Z(n437) );
  XOR2_X1 U488 ( .A(G197GAT), .B(G141GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(G169GAT), .B(G50GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U491 ( .A(KEYINPUT29), .B(G8GAT), .Z(n433) );
  XNOR2_X1 U492 ( .A(G113GAT), .B(G1GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n438), .B(KEYINPUT30), .Z(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT67), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n574) );
  XNOR2_X1 U499 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n453) );
  NAND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n293), .B(n443), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n447) );
  XNOR2_X1 U504 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n446) );
  XOR2_X1 U505 ( .A(n452), .B(n451), .Z(n579) );
  XOR2_X1 U506 ( .A(n453), .B(n579), .Z(n563) );
  INV_X1 U507 ( .A(n563), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n574), .A2(n454), .ZN(n518) );
  XOR2_X1 U509 ( .A(KEYINPUT107), .B(n455), .Z(n537) );
  NAND2_X1 U510 ( .A1(n537), .A2(n526), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(n350), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n458), .B(n457), .ZN(G1339GAT) );
  INV_X1 U514 ( .A(KEYINPUT54), .ZN(n473) );
  XNOR2_X1 U515 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n574), .A2(n563), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n585), .B(KEYINPUT111), .ZN(n570) );
  NOR2_X1 U519 ( .A1(n461), .A2(n570), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT113), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n463), .A2(n556), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT47), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n585), .A2(n589), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n579), .A2(n296), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n574), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n480) );
  INV_X1 U529 ( .A(n471), .ZN(n495) );
  NOR2_X1 U530 ( .A1(n480), .A2(n495), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n573), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n536), .ZN(n562) );
  INV_X1 U535 ( .A(n562), .ZN(n569) );
  NAND2_X1 U536 ( .A1(n556), .A2(n569), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n482), .B(KEYINPUT114), .ZN(n549) );
  AND2_X1 U539 ( .A1(n536), .A2(n549), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT115), .ZN(n484) );
  INV_X1 U541 ( .A(n545), .ZN(n540) );
  NOR2_X1 U542 ( .A1(n540), .A2(n563), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1341GAT) );
  NOR2_X1 U545 ( .A1(n574), .A2(n579), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT72), .B(n488), .Z(n505) );
  NOR2_X1 U547 ( .A1(n585), .A2(n556), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT16), .ZN(n492) );
  INV_X1 U549 ( .A(n490), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n492), .A2(n491), .ZN(n517) );
  NOR2_X1 U551 ( .A1(n505), .A2(n517), .ZN(n500) );
  NAND2_X1 U552 ( .A1(n532), .A2(n500), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  XOR2_X1 U555 ( .A(G8GAT), .B(KEYINPUT95), .Z(n497) );
  NAND2_X1 U556 ( .A1(n500), .A2(n471), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U559 ( .A1(n500), .A2(n536), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n502) );
  NAND2_X1 U562 ( .A1(n500), .A2(n526), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT99), .Z(n508) );
  NOR2_X1 U566 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(KEYINPUT38), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n515), .A2(n532), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U570 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NAND2_X1 U572 ( .A1(n515), .A2(n471), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n513) );
  NAND2_X1 U575 ( .A1(n515), .A2(n536), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(n514), .ZN(G1330GAT) );
  NAND2_X1 U578 ( .A1(n526), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n516), .ZN(G1331GAT) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n527), .A2(n532), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1332GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n522) );
  NAND2_X1 U585 ( .A1(n527), .A2(n471), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G64GAT), .B(n523), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n536), .A2(n527), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT104), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G71GAT), .B(n525), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT105), .Z(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n537), .A2(n532), .ZN(n533) );
  XNOR2_X1 U597 ( .A(KEYINPUT108), .B(n533), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G85GAT), .B(n534), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n471), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U601 ( .A(G99GAT), .B(KEYINPUT109), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1338GAT) );
  NOR2_X1 U604 ( .A1(n574), .A2(n540), .ZN(n541) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n541), .Z(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U607 ( .A1(n545), .A2(n570), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n556), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n572), .ZN(n557) );
  NOR2_X1 U615 ( .A1(n574), .A2(n557), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n563), .A2(n557), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n585), .A2(n557), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  INV_X1 U624 ( .A(n556), .ZN(n558) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT120), .B(n559), .Z(n560) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n574), .A2(n562), .ZN(n561) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT56), .B(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n588) );
  NOR2_X1 U639 ( .A1(n588), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  INV_X1 U644 ( .A(n579), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n588), .A2(n580), .ZN(n584) );
  XOR2_X1 U646 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n588), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(n586), .Z(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

