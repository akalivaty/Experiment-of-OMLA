//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G110), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  XNOR2_X1  g010(.A(G119), .B(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G125), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT77), .A4(G125), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  OAI21_X1  g022(.A(G140), .B1(new_n208), .B2(KEYINPUT76), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n202), .A3(G125), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT16), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(G146), .A3(new_n206), .A4(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n200), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n194), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n217));
  XOR2_X1   g031(.A(G125), .B(G140), .Z(new_n218));
  OR2_X1    g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT78), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n206), .A3(new_n205), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n199), .B1(new_n225), .B2(new_n214), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n217), .A2(new_n214), .A3(new_n219), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT22), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n221), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n216), .A2(new_n220), .A3(new_n232), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n187), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT79), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT25), .B1(new_n241), .B2(KEYINPUT80), .ZN(new_n242));
  OAI22_X1  g056(.A1(new_n239), .A2(new_n240), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n235), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n234), .A2(new_n236), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT81), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n245), .A2(G902), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n253));
  INV_X1    g067(.A(G113), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(KEYINPUT2), .B2(G113), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n255), .A2(new_n257), .B1(KEYINPUT2), .B2(G113), .ZN(new_n258));
  XNOR2_X1  g072(.A(G116), .B(G119), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n258), .A2(new_n259), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(G137), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT11), .A3(G134), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(new_n268), .A3(new_n271), .A4(new_n266), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  XNOR2_X1  g088(.A(G143), .B(G146), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n224), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G146), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT0), .B(G128), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT64), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n262), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n192), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n278), .A3(new_n280), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(KEYINPUT1), .A3(G146), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n264), .A2(G137), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n267), .A2(G134), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n272), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n272), .A2(new_n294), .A3(KEYINPUT68), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n291), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n252), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT72), .B(new_n252), .C1(new_n286), .C2(new_n299), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n273), .A2(new_n284), .A3(KEYINPUT67), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT67), .B1(new_n273), .B2(new_n284), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n272), .A2(new_n294), .A3(KEYINPUT68), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT68), .B1(new_n272), .B2(new_n294), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n307), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n260), .A2(new_n261), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n307), .A2(new_n262), .A3(new_n312), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n304), .B1(new_n319), .B2(KEYINPUT28), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n229), .A3(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G902), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n307), .A2(KEYINPUT30), .A3(new_n312), .A4(new_n314), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n272), .A2(new_n294), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n273), .A2(new_n284), .B1(new_n333), .B2(new_n308), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n334), .B2(KEYINPUT30), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n308), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n285), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT65), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n340), .A3(new_n316), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n318), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n327), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n316), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n318), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT28), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n302), .A2(new_n303), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n326), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n328), .B(new_n343), .C1(new_n348), .C2(KEYINPUT75), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n330), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G472), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n252), .B1(new_n318), .B2(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n327), .B1(new_n353), .B2(new_n304), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT73), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT73), .B(new_n327), .C1(new_n353), .C2(new_n304), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n318), .A2(new_n326), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT31), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n341), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n341), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT31), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G472), .A2(G902), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n352), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n251), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n213), .A2(new_n215), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n322), .A2(new_n229), .A3(G214), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G143), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(new_n271), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n271), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n376), .B(new_n380), .C1(new_n381), .C2(KEYINPUT17), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n209), .A2(new_n211), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n219), .B1(new_n388), .B2(new_n224), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n386), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n382), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n214), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT19), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n218), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(KEYINPUT19), .B2(new_n388), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G146), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n391), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n385), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n381), .B(new_n214), .C1(G146), .C2(new_n396), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n391), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(G475), .A2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT20), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n391), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT94), .B1(new_n401), .B2(new_n391), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(new_n385), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n407), .B(new_n404), .C1(new_n410), .C2(new_n392), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G475), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n385), .B1(new_n382), .B2(new_n391), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n392), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n415), .B2(new_n235), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n419), .A2(G952), .A3(new_n229), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT9), .B(G234), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT82), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G217), .A3(new_n229), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT99), .ZN(new_n428));
  INV_X1    g242(.A(G116), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G122), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n430), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G107), .B1(new_n430), .B2(new_n435), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT97), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n431), .A2(G116), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n433), .B1(new_n440), .B2(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n430), .A2(new_n432), .A3(new_n435), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n434), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n192), .A2(G143), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n279), .A2(KEYINPUT95), .A3(G128), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT95), .B1(new_n279), .B2(G128), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G134), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n192), .B2(G143), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n279), .A2(KEYINPUT95), .A3(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n264), .A3(new_n445), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT98), .B1(new_n444), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n434), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT97), .B1(new_n436), .B2(new_n437), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(new_n439), .A3(new_n442), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT98), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n454), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n430), .A2(new_n432), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n434), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT13), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT96), .B1(new_n453), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n469), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT96), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n451), .A2(new_n452), .A3(new_n472), .A4(KEYINPUT13), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n445), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n468), .B1(new_n474), .B2(G134), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n428), .B1(new_n464), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT99), .B(new_n475), .C1(new_n456), .C2(new_n463), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n427), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n458), .A2(new_n459), .ZN(new_n480));
  AND4_X1   g294(.A1(new_n461), .A2(new_n480), .A3(new_n462), .A4(new_n434), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT99), .ZN(new_n484));
  INV_X1    g298(.A(new_n427), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n235), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT102), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n464), .A2(new_n428), .A3(new_n476), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n485), .B1(new_n484), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n477), .A2(new_n427), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n235), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT100), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT100), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n235), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n493), .B1(new_n501), .B2(new_n489), .ZN(new_n502));
  AOI211_X1 g316(.A(KEYINPUT101), .B(new_n490), .C1(new_n498), .C2(new_n500), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n424), .B(new_n492), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G210), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n258), .A2(new_n259), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n429), .A2(KEYINPUT5), .A3(G119), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n254), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(KEYINPUT84), .A2(G101), .ZN(new_n514));
  NOR2_X1   g328(.A1(KEYINPUT84), .A2(G101), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT3), .B1(new_n384), .B2(G107), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n384), .A2(G107), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT3), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n433), .A3(G104), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n433), .A2(G104), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n524), .B2(G101), .ZN(new_n525));
  INV_X1    g339(.A(G101), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT85), .B(new_n526), .C1(new_n523), .C2(new_n518), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT86), .B(new_n521), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G104), .B(G107), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT85), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n522), .A3(G101), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT86), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n513), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n517), .A2(new_n520), .A3(new_n518), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G101), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT4), .A3(new_n521), .ZN(new_n538));
  OAI221_X1 g352(.A(new_n538), .B1(KEYINPUT4), .B2(new_n537), .C1(new_n261), .C2(new_n260), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G110), .B(G122), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT90), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n535), .A2(new_n539), .A3(new_n541), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n277), .A2(new_n283), .A3(G125), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(G125), .B2(new_n308), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT91), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n229), .A2(G224), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT92), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n546), .A2(new_n547), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n550), .A2(KEYINPUT7), .A3(new_n552), .A4(new_n554), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n549), .B1(new_n561), .B2(new_n557), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n508), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n259), .A2(KEYINPUT93), .A3(KEYINPUT5), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n510), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n507), .B(new_n567), .C1(new_n529), .C2(new_n534), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n533), .A2(new_n521), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n512), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n541), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n535), .A2(new_n539), .A3(new_n541), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n235), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n506), .B1(new_n559), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n558), .A2(new_n555), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n574), .A2(KEYINPUT6), .B1(new_n540), .B2(new_n542), .ZN(new_n579));
  INV_X1    g393(.A(new_n547), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n572), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n568), .B2(new_n570), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n544), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n584), .B2(new_n563), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n585), .A3(new_n505), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G214), .B1(G237), .B2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n504), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n426), .A2(new_n235), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n591), .A2(G221), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n229), .A2(G227), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G140), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT83), .B(G110), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n529), .A2(new_n534), .A3(new_n308), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n533), .A2(new_n308), .A3(new_n521), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n273), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n569), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n291), .A3(new_n528), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n599), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT12), .A3(new_n273), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT10), .B(new_n308), .C1(new_n529), .C2(new_n534), .ZN(new_n610));
  INV_X1    g424(.A(new_n273), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n536), .A2(G101), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT4), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n612), .A2(new_n613), .B1(new_n283), .B2(new_n277), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n538), .A2(new_n614), .B1(new_n599), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT87), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n610), .A2(new_n616), .A3(new_n619), .A4(new_n611), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n609), .A2(KEYINPUT88), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT88), .B1(new_n609), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n597), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n597), .B1(new_n618), .B2(new_n620), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n610), .A2(new_n616), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n273), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(G469), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT89), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n597), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT88), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n618), .A2(new_n620), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT12), .B1(new_n607), .B2(new_n273), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n602), .B(new_n611), .C1(new_n606), .C2(new_n599), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n609), .A2(new_n621), .A3(KEYINPUT88), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n628), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n235), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT89), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(G469), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n625), .A2(new_n609), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n632), .B1(new_n621), .B2(new_n627), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n630), .B(new_n235), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n631), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n375), .A2(new_n590), .A3(new_n593), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(new_n516), .Z(G3));
  INV_X1    g464(.A(new_n647), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n642), .A2(G469), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(KEYINPUT89), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n592), .B1(new_n653), .B2(new_n644), .ZN(new_n654));
  AOI21_X1  g468(.A(G478), .B1(new_n498), .B2(new_n500), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n488), .A2(G902), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n427), .A2(KEYINPUT104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n483), .B(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n479), .A2(new_n660), .A3(new_n486), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n418), .B1(new_n655), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n588), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n505), .B1(new_n581), .B2(new_n585), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(KEYINPUT103), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n577), .A2(new_n669), .A3(new_n586), .ZN(new_n670));
  INV_X1    g484(.A(new_n423), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n367), .B2(new_n235), .ZN(new_n675));
  INV_X1    g489(.A(new_n368), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n360), .B1(new_n359), .B2(new_n341), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(KEYINPUT71), .B2(new_n361), .ZN(new_n678));
  INV_X1    g492(.A(new_n366), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n676), .B1(new_n680), .B2(new_n358), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n675), .A2(new_n681), .A3(new_n251), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n654), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n491), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n499), .B1(new_n487), .B2(new_n235), .ZN(new_n688));
  AOI211_X1 g502(.A(KEYINPUT100), .B(G902), .C1(new_n479), .C2(new_n486), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n489), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n501), .A2(new_n493), .A3(new_n489), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n418), .A3(new_n672), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n654), .A2(new_n682), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT35), .B(G107), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G9));
  NAND2_X1  g511(.A1(new_n221), .A2(new_n228), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n249), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n246), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n675), .A2(new_n681), .A3(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n590), .A2(new_n593), .A3(new_n648), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n352), .B(new_n369), .C1(new_n681), .C2(new_n372), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n702), .A2(new_n668), .A3(new_n670), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n648), .A2(new_n709), .A3(new_n593), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n416), .B1(new_n406), .B2(new_n411), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n420), .B1(new_n421), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n708), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n693), .A2(new_n418), .A3(new_n716), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n710), .B1(new_n370), .B2(new_n374), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G128), .ZN(G30));
  XOR2_X1   g538(.A(new_n716), .B(KEYINPUT39), .Z(new_n725));
  NAND2_X1  g539(.A1(new_n654), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT40), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n319), .A2(new_n327), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n363), .A3(G472), .ZN(new_n729));
  NAND2_X1  g543(.A1(G472), .A2(G902), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT106), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(new_n369), .C1(new_n681), .C2(new_n372), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT107), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n587), .B(KEYINPUT38), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n588), .A3(new_n703), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n734), .A2(new_n693), .A3(new_n714), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n727), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G143), .ZN(G45));
  OAI211_X1 g553(.A(new_n418), .B(new_n717), .C1(new_n655), .C2(new_n664), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n712), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n224), .ZN(G48));
  INV_X1    g556(.A(new_n251), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n621), .A2(new_n627), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n744), .A2(new_n597), .B1(new_n625), .B2(new_n609), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n745), .B2(G902), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n593), .A3(new_n647), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n709), .A2(new_n673), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND3_X1  g565(.A1(new_n694), .A2(new_n375), .A3(new_n748), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NOR2_X1   g567(.A1(new_n710), .A2(new_n747), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n709), .A2(new_n754), .A3(new_n693), .A4(new_n424), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  INV_X1    g570(.A(new_n504), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n709), .A4(new_n754), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  NOR2_X1   g575(.A1(new_n747), .A2(new_n423), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n668), .A2(new_n670), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n713), .A2(new_n762), .A3(new_n418), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n675), .A2(new_n251), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n364), .A2(new_n361), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n320), .A2(new_n326), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n368), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n431), .ZN(G24));
  NOR3_X1   g586(.A1(new_n740), .A2(new_n763), .A3(new_n747), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n702), .A2(new_n769), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n675), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT109), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n740), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n747), .A2(new_n763), .ZN(new_n778));
  AND4_X1   g592(.A1(KEYINPUT109), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n208), .ZN(G27));
  AOI21_X1  g595(.A(new_n651), .B1(new_n642), .B2(G469), .ZN(new_n782));
  INV_X1    g596(.A(new_n587), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n592), .A2(new_n666), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n709), .A3(new_n743), .A4(new_n777), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n782), .A2(new_n740), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n371), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n251), .B1(new_n370), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n271), .ZN(G33));
  AND3_X1   g608(.A1(new_n720), .A2(new_n375), .A3(new_n786), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n264), .ZN(G36));
  NAND2_X1  g610(.A1(new_n783), .A2(new_n588), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n675), .A2(new_n681), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n702), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT112), .Z(new_n800));
  OAI21_X1  g614(.A(new_n488), .B1(new_n688), .B2(new_n689), .ZN(new_n801));
  INV_X1    g615(.A(new_n663), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n656), .B1(new_n802), .B2(new_n661), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n714), .ZN(new_n805));
  NAND2_X1  g619(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n800), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n797), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n640), .B2(new_n641), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n624), .A2(KEYINPUT45), .A3(new_n628), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(G469), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(G469), .A2(G902), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n651), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n817), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n592), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n725), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n800), .A2(KEYINPUT44), .A3(new_n809), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n812), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT113), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(new_n267), .ZN(G39));
  OR2_X1    g643(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n830));
  NAND2_X1  g644(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n822), .A2(new_n831), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n709), .A2(new_n743), .A3(new_n740), .A4(new_n797), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n838));
  INV_X1    g652(.A(new_n780), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n652), .A2(new_n647), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n702), .A2(new_n592), .A3(new_n716), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n733), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n713), .A2(new_n418), .A3(new_n764), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n712), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n777), .ZN(new_n846));
  AND4_X1   g660(.A1(KEYINPUT52), .A2(new_n723), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n848));
  AOI21_X1  g662(.A(new_n780), .B1(new_n719), .B2(new_n722), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n846), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n649), .A2(new_n705), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n665), .B1(new_n693), .B2(new_n418), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n589), .A2(new_n423), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n648), .A2(new_n593), .A3(new_n682), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT116), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n654), .B(new_n590), .C1(new_n375), .C2(new_n704), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n654), .A2(new_n682), .A3(new_n853), .A4(new_n854), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n749), .B1(new_n765), .B2(new_n770), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(new_n760), .A3(new_n752), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n786), .A2(new_n777), .A3(new_n775), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n797), .A2(new_n418), .A3(new_n716), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n709), .A3(new_n693), .A4(new_n702), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n648), .A2(new_n593), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n793), .A2(new_n795), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n866), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n838), .B1(new_n851), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n859), .A2(new_n861), .A3(new_n860), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n861), .B1(new_n859), .B2(new_n860), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n872), .B(new_n866), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n723), .A2(new_n839), .A3(new_n846), .ZN(new_n879));
  INV_X1    g693(.A(new_n848), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n846), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n883), .A3(KEYINPUT120), .A4(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n863), .A2(KEYINPUT117), .A3(new_n866), .A4(new_n872), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n882), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n887), .A2(new_n888), .A3(new_n883), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n893), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n893), .B2(new_n892), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT119), .B1(new_n898), .B2(new_n893), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n809), .A2(new_n420), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n904), .A2(new_n766), .A3(new_n769), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n735), .A2(new_n588), .A3(new_n747), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT50), .Z(new_n908));
  NOR2_X1   g722(.A1(new_n797), .A2(new_n747), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n734), .A2(new_n743), .A3(new_n420), .A4(new_n909), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n910), .A2(new_n418), .A3(new_n804), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n904), .A2(new_n775), .A3(new_n909), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n746), .A2(new_n647), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT115), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n834), .B1(new_n592), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n905), .A2(new_n588), .A3(new_n783), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n913), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n913), .B2(new_n919), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n904), .A2(new_n792), .A3(new_n909), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT48), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n905), .A2(new_n778), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(G952), .A3(new_n229), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n910), .A2(new_n665), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n903), .A2(new_n929), .B1(G952), .B2(G953), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n915), .B(KEYINPUT49), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n743), .A2(new_n784), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(new_n735), .A3(new_n805), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n734), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G75));
  NOR2_X1   g749(.A1(new_n229), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n874), .A2(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n938));
  INV_X1    g752(.A(G210), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n235), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n579), .A2(new_n580), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n578), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT56), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT56), .B1(new_n940), .B2(KEYINPUT121), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n895), .A2(G902), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n950), .B2(new_n943), .ZN(G51));
  XNOR2_X1  g765(.A(new_n938), .B(KEYINPUT54), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n817), .B(KEYINPUT57), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n952), .A2(new_n953), .B1(new_n646), .B2(new_n645), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n948), .A2(new_n816), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n936), .B1(new_n954), .B2(new_n955), .ZN(G54));
  INV_X1    g770(.A(new_n948), .ZN(new_n957));
  INV_X1    g771(.A(new_n403), .ZN(new_n958));
  AND2_X1   g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n936), .ZN(G60));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n802), .B2(new_n661), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n937), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n903), .A2(new_n965), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n802), .A2(new_n661), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G63));
  XNOR2_X1  g784(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n244), .A2(new_n235), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n895), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n936), .B1(new_n974), .B2(new_n248), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n885), .B2(new_n894), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT123), .B1(new_n977), .B2(new_n700), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n979));
  INV_X1    g793(.A(new_n700), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n938), .A2(new_n979), .A3(new_n980), .A4(new_n976), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n975), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n975), .B(KEYINPUT61), .C1(new_n978), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  NAND2_X1  g800(.A1(new_n863), .A2(new_n866), .ZN(new_n987));
  NAND2_X1  g801(.A1(G224), .A2(G953), .ZN(new_n988));
  OAI22_X1  g802(.A1(new_n987), .A2(G953), .B1(new_n422), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n941), .B1(G898), .B2(new_n229), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(G69));
  AOI211_X1 g805(.A(new_n741), .B(new_n780), .C1(new_n719), .C2(new_n722), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n738), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n375), .A2(new_n853), .A3(new_n588), .A4(new_n783), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(new_n726), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n834), .B2(new_n835), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n994), .A2(new_n827), .A3(new_n995), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n229), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n331), .A2(new_n340), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n396), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n229), .A2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n843), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n825), .A2(new_n1006), .A3(new_n792), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n793), .A2(new_n795), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n834), .B2(new_n835), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n827), .A2(new_n1007), .A3(new_n992), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1005), .B1(new_n1010), .B2(new_n229), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(new_n1002), .A3(new_n1013), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1022), .A2(KEYINPUT125), .A3(new_n1017), .A4(new_n1004), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1020), .A2(new_n1023), .ZN(G72));
  XOR2_X1   g838(.A(new_n730), .B(KEYINPUT63), .Z(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n999), .B2(new_n987), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n342), .B(KEYINPUT126), .Z(new_n1027));
  NAND3_X1  g841(.A1(new_n1026), .A2(new_n326), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1025), .B1(new_n1010), .B2(new_n987), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1027), .A2(new_n326), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n936), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n900), .A2(new_n901), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1025), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n343), .A2(KEYINPUT127), .ZN(new_n1035));
  AOI22_X1  g849(.A1(new_n343), .A2(KEYINPUT127), .B1(new_n341), .B2(new_n359), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1032), .B1(new_n1033), .B2(new_n1037), .ZN(G57));
endmodule


