//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n195), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G134), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n203), .A2(new_n204), .A3(new_n197), .A4(new_n196), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n212), .A2(new_n214), .B1(new_n208), .B2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(new_n207), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n210), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n206), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G146), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n211), .A2(G143), .ZN(new_n222));
  OAI211_X1 g036(.A(G128), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n212), .B(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n201), .A2(new_n197), .A3(KEYINPUT66), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n195), .A3(G134), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(G131), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n205), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G116), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G119), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G113), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n233), .B(new_n235), .C1(new_n237), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n233), .A2(new_n235), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n219), .A2(new_n231), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n217), .A2(new_n216), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n221), .B2(new_n222), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n251), .B2(new_n209), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n199), .B2(new_n205), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n205), .A2(new_n225), .A3(new_n223), .A4(new_n230), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n244), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n247), .B1(new_n255), .B2(new_n246), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n248), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI211_X1 g078(.A(KEYINPUT68), .B(new_n247), .C1(new_n255), .C2(new_n246), .ZN(new_n265));
  OR4_X1    g079(.A1(KEYINPUT70), .A2(new_n258), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n255), .A2(new_n246), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  INV_X1    g083(.A(new_n265), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n263), .A3(new_n270), .A4(new_n248), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT30), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n219), .B2(new_n231), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n244), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n246), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n264), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n266), .A2(new_n272), .A3(new_n273), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n246), .A2(new_n281), .A3(new_n247), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n268), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n284), .A2(new_n273), .A3(new_n264), .ZN(new_n285));
  XOR2_X1   g099(.A(KEYINPUT72), .B(G902), .Z(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n187), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n264), .B1(new_n258), .B2(new_n265), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n246), .A2(new_n292), .A3(new_n263), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT30), .B1(new_n253), .B2(new_n254), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n219), .A2(new_n231), .A3(new_n275), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n245), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n246), .A2(new_n263), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT31), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n246), .A2(new_n292), .A3(new_n263), .ZN(new_n301));
  AND4_X1   g115(.A1(KEYINPUT31), .A2(new_n277), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n291), .B(KEYINPUT69), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n277), .A2(new_n299), .A3(new_n301), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n277), .A2(new_n299), .A3(KEYINPUT31), .A4(new_n301), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT69), .B1(new_n309), .B2(new_n291), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n290), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT32), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n291), .B1(new_n300), .B2(new_n302), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n303), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT32), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n290), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n289), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G217), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n286), .B2(G234), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(new_n211), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n232), .B2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n330), .B(new_n331), .C1(G119), .C2(new_n224), .ZN(new_n332));
  XNOR2_X1  g146(.A(G119), .B(G128), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  OAI22_X1  g148(.A1(new_n332), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT16), .B1(new_n322), .B2(G125), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n324), .B2(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n322), .A2(KEYINPUT73), .A3(G125), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n325), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(new_n211), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n342), .B(new_n211), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n332), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT74), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI211_X1 g162(.A(G146), .B(new_n337), .C1(new_n341), .C2(KEYINPUT16), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT74), .B(new_n347), .C1(new_n343), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n353), .B(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n347), .B1(new_n343), .B2(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n350), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n345), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT25), .B1(new_n366), .B2(new_n286), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n363), .B2(new_n345), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n344), .B(new_n358), .C1(new_n362), .C2(new_n350), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT25), .B(new_n286), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n321), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n321), .A2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  INV_X1    g190(.A(G237), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n354), .A3(G214), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n213), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT18), .A3(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n326), .B(KEYINPUT75), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n341), .A2(G146), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n382), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n341), .A2(KEYINPUT19), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT19), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n323), .A2(new_n325), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n211), .A3(new_n390), .ZN(new_n391));
  AND4_X1   g205(.A1(G143), .A2(new_n377), .A3(new_n354), .A4(G214), .ZN(new_n392));
  AOI21_X1  g206(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n393));
  OAI21_X1  g207(.A(G131), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n379), .A2(new_n204), .A3(new_n380), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n391), .B(new_n396), .C1(new_n211), .C2(new_n342), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT17), .B(G131), .C1(new_n392), .C2(new_n393), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT87), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n394), .A2(new_n406), .A3(new_n395), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n383), .A2(new_n408), .A3(KEYINPUT17), .A4(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n401), .B(new_n387), .C1(new_n346), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n376), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT20), .B(new_n415), .C1(new_n403), .C2(new_n411), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n387), .B1(new_n346), .B2(new_n410), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n402), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n414), .A2(new_n416), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT88), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n423), .B1(new_n420), .B2(new_n417), .C1(new_n414), .C2(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G128), .B(G143), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(new_n189), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n234), .A2(KEYINPUT14), .A3(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(G116), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(G107), .B(new_n428), .C1(new_n430), .C2(KEYINPUT14), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n427), .B(new_n431), .C1(G107), .C2(new_n430), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(G128), .A3(new_n213), .ZN(new_n434));
  INV_X1    g248(.A(new_n426), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n434), .B(G134), .C1(new_n435), .C2(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n189), .ZN(new_n437));
  INV_X1    g251(.A(G107), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n429), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT9), .B(G234), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(new_n320), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n432), .A2(new_n440), .A3(new_n443), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n287), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G478), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT15), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n447), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G234), .A2(G237), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(G952), .A3(new_n354), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n287), .A2(G953), .A3(new_n452), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT90), .Z(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(G898), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n425), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT5), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(G113), .C1(KEYINPUT5), .C2(new_n233), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n400), .A2(G107), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n400), .A2(G107), .ZN(new_n467));
  OAI21_X1  g281(.A(G101), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT79), .B(G101), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT3), .B1(new_n400), .B2(G107), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n438), .A3(G104), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n469), .A2(new_n465), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n464), .A2(new_n240), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n464), .A2(new_n240), .B1(new_n473), .B2(new_n468), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n249), .B(G125), .C1(new_n251), .C2(new_n209), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n223), .A2(new_n225), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(G125), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G224), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(KEYINPUT7), .C1(new_n481), .C2(G953), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n470), .A2(new_n472), .A3(new_n465), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G101), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n473), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n487), .A3(G101), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n244), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n474), .B(new_n460), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n477), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n481), .A2(G953), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n493));
  OAI221_X1 g307(.A(new_n478), .B1(new_n492), .B2(new_n493), .C1(G125), .C2(new_n479), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G210), .B1(G237), .B2(G902), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n474), .B1(new_n486), .B2(new_n489), .ZN(new_n499));
  INV_X1    g313(.A(new_n460), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n480), .B(new_n492), .Z(new_n503));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n497), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n498), .B1(new_n497), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G214), .B1(G237), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G221), .B1(new_n442), .B2(G902), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT78), .Z(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G140), .ZN(new_n515));
  INV_X1    g329(.A(G227), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G953), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n515), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n473), .A2(new_n468), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n479), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n473), .A2(new_n468), .A3(new_n223), .A4(new_n225), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n206), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n522), .A2(KEYINPUT82), .A3(new_n524), .A4(new_n206), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n531));
  NAND2_X1  g345(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT81), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n485), .A2(new_n218), .A3(new_n488), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n468), .A4(new_n473), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n206), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n518), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n206), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n536), .A2(new_n537), .ZN(new_n542));
  INV_X1    g356(.A(new_n206), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n533), .A4(new_n535), .ZN(new_n544));
  INV_X1    g358(.A(new_n518), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(G469), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  INV_X1    g362(.A(G902), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n527), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n525), .B(new_n553), .C1(new_n522), .C2(new_n206), .ZN(new_n554));
  INV_X1    g368(.A(new_n529), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT83), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n528), .A2(new_n557), .A3(new_n529), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n556), .A2(new_n544), .A3(new_n545), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n541), .A2(new_n544), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n518), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n548), .A3(new_n286), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n514), .B1(new_n552), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n459), .A2(new_n512), .A3(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n319), .A2(new_n375), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT91), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(new_n469), .ZN(G3));
  OAI21_X1  g382(.A(new_n286), .B1(new_n304), .B2(new_n310), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n569), .A2(G472), .B1(new_n316), .B2(new_n290), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n564), .A2(new_n374), .A3(new_n372), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT92), .Z(new_n573));
  INV_X1    g387(.A(new_n457), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n287), .A2(new_n448), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n445), .A2(new_n576), .A3(new_n446), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n445), .B2(new_n446), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n580));
  INV_X1    g394(.A(new_n447), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n448), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n447), .A2(KEYINPUT94), .A3(G478), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n422), .A2(new_n424), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n497), .A2(new_n506), .A3(new_n498), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n510), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n509), .B2(new_n588), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n573), .A2(new_n574), .A3(new_n586), .A4(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT34), .B(G104), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G6));
  INV_X1    g407(.A(new_n414), .ZN(new_n594));
  INV_X1    g408(.A(new_n416), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n420), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G475), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n596), .A2(new_n598), .A3(new_n574), .A4(new_n451), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n421), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n602), .A2(KEYINPUT95), .A3(new_n574), .A4(new_n451), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n573), .A2(new_n590), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G107), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  NOR2_X1   g421(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n352), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n373), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n372), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n287), .B1(new_n315), .B2(new_n303), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n311), .B(new_n611), .C1(new_n612), .C2(new_n187), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n565), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT37), .B(G110), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  NAND2_X1  g432(.A1(new_n280), .A2(new_n288), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n317), .B1(new_n316), .B2(new_n290), .ZN(new_n621));
  INV_X1    g435(.A(new_n290), .ZN(new_n622));
  AOI211_X1 g436(.A(KEYINPUT32), .B(new_n622), .C1(new_n315), .C2(new_n303), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n453), .B(KEYINPUT96), .Z(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n455), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n602), .A2(new_n451), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n564), .A2(new_n611), .A3(new_n590), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  AOI22_X1  g448(.A1(new_n297), .A2(new_n299), .B1(new_n264), .B2(new_n267), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n636), .B1(new_n621), .B2(new_n623), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n628), .B(KEYINPUT39), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n564), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT40), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n422), .A2(new_n424), .A3(new_n451), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n611), .A2(new_n511), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n497), .A2(new_n506), .ZN(new_n644));
  INV_X1    g458(.A(new_n498), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n587), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n638), .A2(new_n641), .A3(new_n642), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n213), .ZN(G45));
  AND4_X1   g465(.A1(new_n422), .A2(new_n424), .A3(new_n584), .A4(new_n629), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n564), .A3(new_n611), .A4(new_n590), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n624), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  NAND2_X1  g470(.A1(new_n312), .A2(new_n318), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n375), .B1(new_n657), .B2(new_n620), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n548), .B1(new_n562), .B2(new_n286), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n513), .A3(new_n563), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n510), .B(new_n662), .C1(new_n647), .C2(KEYINPUT93), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n661), .A2(new_n663), .A3(new_n585), .A4(new_n457), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT41), .B(G113), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT97), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G15));
  AOI211_X1 g482(.A(G469), .B(new_n287), .C1(new_n559), .C2(new_n561), .ZN(new_n669));
  INV_X1    g483(.A(new_n513), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n659), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n604), .A2(new_n671), .A3(new_n590), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT98), .B(G116), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G18));
  AND4_X1   g489(.A1(new_n459), .A2(new_n671), .A3(new_n590), .A4(new_n611), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n624), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  OAI21_X1  g492(.A(KEYINPUT100), .B1(new_n663), .B2(new_n642), .ZN(new_n679));
  INV_X1    g493(.A(new_n425), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n590), .A3(new_n681), .A4(new_n451), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n375), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n300), .A2(new_n302), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n284), .A2(new_n264), .ZN(new_n686));
  OAI211_X1 g500(.A(KEYINPUT99), .B(new_n290), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT99), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n307), .A2(new_n308), .B1(new_n264), .B2(new_n284), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n622), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(G472), .B2(new_n569), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n661), .A2(new_n457), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n683), .A2(new_n684), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  NOR2_X1   g509(.A1(new_n661), .A2(new_n663), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n692), .A2(new_n696), .A3(new_n611), .A4(new_n652), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  NAND2_X1  g512(.A1(new_n540), .A2(new_n546), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n546), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(G469), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n563), .A3(new_n551), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n509), .A2(new_n705), .A3(new_n510), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT102), .B1(new_n647), .B2(new_n511), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n513), .A2(new_n704), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n624), .A2(new_n684), .A3(new_n708), .A4(new_n652), .ZN(new_n709));
  NOR2_X1   g523(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n710), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n658), .A2(new_n652), .A3(new_n712), .A4(new_n708), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n711), .A2(new_n713), .A3(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  AND4_X1   g533(.A1(new_n684), .A2(new_n624), .A3(new_n630), .A4(new_n708), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n189), .ZN(G36));
  INV_X1    g535(.A(new_n570), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n425), .A2(KEYINPUT105), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n422), .B2(new_n424), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n584), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT43), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n425), .A2(new_n728), .A3(new_n584), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n722), .A2(new_n727), .A3(new_n611), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n702), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n548), .B1(new_n699), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n550), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n563), .B1(new_n736), .B2(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n513), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n707), .A2(new_n706), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n740), .A2(new_n639), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n731), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT106), .B(G137), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G39));
  NAND4_X1  g560(.A1(new_n319), .A2(new_n375), .A3(new_n652), .A4(new_n742), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n755));
  NOR2_X1   g569(.A1(G952), .A2(G953), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n711), .A2(new_n713), .A3(KEYINPUT104), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT104), .B1(new_n711), .B2(new_n713), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n647), .A2(new_n574), .A3(new_n510), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n586), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT109), .B1(new_n761), .B2(new_n585), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n570), .A2(new_n571), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n760), .B1(new_n566), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n624), .A2(new_n615), .A3(new_n684), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n570), .A2(new_n571), .A3(new_n764), .A4(new_n765), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n624), .B(new_n684), .C1(new_n664), .C2(new_n672), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n694), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n425), .A2(new_n451), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n570), .A2(new_n571), .A3(new_n762), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n677), .A2(new_n616), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n569), .A2(G472), .ZN(new_n778));
  INV_X1    g592(.A(new_n691), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n611), .A4(new_n652), .ZN(new_n780));
  INV_X1    g594(.A(new_n708), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n421), .A2(new_n451), .A3(new_n628), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n742), .A2(new_n564), .A3(new_n611), .A4(new_n782), .ZN(new_n783));
  OAI22_X1  g597(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n319), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n720), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n771), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT111), .B1(new_n759), .B2(new_n786), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n676), .A2(new_n624), .B1(new_n614), .B2(new_n615), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n772), .A3(new_n694), .A4(new_n775), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n767), .B2(new_n770), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n718), .A2(new_n790), .A3(new_n791), .A4(new_n785), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n704), .A2(new_n513), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n611), .B2(new_n628), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n372), .A2(KEYINPUT112), .A3(new_n610), .A4(new_n629), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n637), .A2(new_n683), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n624), .B1(new_n632), .B2(new_n654), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n697), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n696), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n780), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n657), .A2(new_n620), .B1(new_n631), .B2(new_n653), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(KEYINPUT52), .A3(new_n798), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(new_n806), .B2(new_n798), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n787), .A2(new_n792), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n771), .A2(new_n777), .A3(new_n785), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n802), .A2(new_n807), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n718), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT114), .A4(KEYINPUT54), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n810), .B1(new_n711), .B2(new_n713), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n815), .A2(new_n812), .A3(new_n809), .A4(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(KEYINPUT52), .A2(new_n798), .A3(new_n799), .A4(new_n697), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n759), .A2(new_n786), .A3(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n821), .B(new_n823), .C1(new_n826), .C2(KEYINPUT53), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n819), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n741), .A2(new_n661), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n727), .A2(new_n626), .A3(new_n729), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n727), .A2(KEYINPUT115), .A3(new_n626), .A4(new_n729), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n658), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT48), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n831), .A2(new_n684), .A3(new_n453), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n638), .A3(new_n586), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(G952), .A3(new_n354), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n692), .A2(new_n684), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n835), .B2(new_n836), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n844), .B2(new_n696), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n692), .A2(new_n611), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n840), .A2(new_n638), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n680), .A2(new_n584), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n837), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n835), .A2(new_n836), .ZN(new_n854));
  INV_X1    g668(.A(new_n843), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n648), .A2(new_n661), .A3(new_n510), .ZN(new_n856));
  AND4_X1   g670(.A1(KEYINPUT50), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT50), .B1(new_n844), .B2(new_n856), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n843), .B(new_n741), .C1(new_n835), .C2(new_n836), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n659), .A2(new_n669), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n514), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n749), .A2(new_n751), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n859), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n868), .B(new_n853), .C1(new_n857), .C2(new_n858), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n863), .B(KEYINPUT116), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n749), .A2(new_n751), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n861), .B2(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n870), .A2(new_n844), .A3(new_n872), .A4(new_n742), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n849), .B(new_n866), .C1(new_n876), .C2(new_n860), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n756), .B1(new_n830), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n375), .A2(new_n511), .A3(new_n514), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT108), .Z(new_n880));
  INV_X1    g694(.A(KEYINPUT49), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n862), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n659), .A2(new_n669), .A3(KEYINPUT49), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n648), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n726), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n884), .A3(new_n638), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n755), .B1(new_n878), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n876), .A2(new_n860), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n866), .A2(new_n849), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n828), .A3(new_n827), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(new_n819), .ZN(new_n894));
  OAI211_X1 g708(.A(KEYINPUT120), .B(new_n886), .C1(new_n894), .C2(new_n756), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n888), .A2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n354), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n817), .A2(new_n810), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n286), .B1(new_n899), .B2(new_n823), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(new_n645), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n502), .A2(new_n505), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n503), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(G51));
  XNOR2_X1  g720(.A(new_n550), .B(KEYINPUT57), .ZN(new_n907));
  INV_X1    g721(.A(new_n827), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n821), .B1(new_n899), .B2(new_n823), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n562), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n900), .A2(new_n733), .A3(new_n735), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(G54));
  AND2_X1   g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n900), .A2(new_n412), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n412), .B1(new_n900), .B2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n897), .ZN(G60));
  OR2_X1    g731(.A1(new_n577), .A2(new_n578), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n908), .B2(new_n909), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n898), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n830), .B2(new_n921), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n927), .A3(new_n898), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(G63));
  XNOR2_X1  g743(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n320), .A2(new_n549), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n899), .B2(new_n823), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n366), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n897), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n934), .A2(KEYINPUT123), .A3(new_n609), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT123), .B1(new_n934), .B2(new_n609), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n936), .B(KEYINPUT61), .C1(new_n938), .C2(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  INV_X1    g757(.A(new_n456), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n354), .B1(new_n944), .B2(G224), .ZN(new_n945));
  INV_X1    g759(.A(new_n790), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n354), .ZN(new_n947));
  INV_X1    g761(.A(G898), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n902), .B1(new_n948), .B2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  NOR2_X1   g764(.A1(new_n274), .A2(new_n276), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n388), .A2(new_n390), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G900), .A2(G953), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n658), .A2(new_n740), .A3(new_n639), .A4(new_n683), .ZN(new_n955));
  INV_X1    g769(.A(new_n806), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n720), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n718), .A2(new_n957), .A3(new_n744), .A4(new_n753), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n953), .B(new_n954), .C1(new_n958), .C2(G953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n650), .A2(new_n956), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n640), .A2(new_n741), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n658), .B(new_n962), .C1(new_n586), .C2(new_n774), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n744), .A2(new_n753), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n959), .B1(new_n967), .B2(new_n953), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT125), .B1(new_n967), .B2(new_n953), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n516), .B2(new_n627), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  OAI221_X1 g787(.A(new_n959), .B1(KEYINPUT125), .B2(new_n971), .C1(new_n967), .C2(new_n953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G72));
  XNOR2_X1  g789(.A(new_n278), .B(KEYINPUT127), .ZN(new_n976));
  OR3_X1    g790(.A1(new_n964), .A2(new_n946), .A3(new_n965), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AND3_X1   g794(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n263), .B(new_n976), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n279), .A2(new_n305), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n814), .A2(new_n818), .A3(new_n980), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n958), .B2(new_n946), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n976), .A2(new_n263), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n897), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(G57));
endmodule


