//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT81), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g010(.A(new_n208), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT80), .B(KEYINPUT2), .Z(new_n213));
  OAI211_X1 g012(.A(new_n203), .B(new_n206), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(G197gat), .ZN(new_n219));
  INV_X1    g018(.A(G204gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G197gat), .A2(G204gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT22), .ZN(new_n223));
  NAND2_X1  g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n224), .ZN(new_n228));
  NOR2_X1   g027(.A1(G211gat), .A2(G218gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n227), .A2(new_n231), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n218), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n225), .A2(new_n226), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n230), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT74), .A3(new_n232), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G228gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n230), .A2(KEYINPUT85), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT85), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n225), .A3(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(new_n216), .C1(new_n225), .C2(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n211), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n210), .A2(new_n214), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n235), .A2(KEYINPUT75), .A3(new_n238), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT75), .B1(new_n235), .B2(new_n238), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n217), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n216), .A3(new_n232), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT3), .B1(new_n257), .B2(KEYINPUT86), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(KEYINPUT86), .B2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n250), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n202), .B(new_n252), .C1(new_n261), .C2(new_n244), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n244), .B1(new_n256), .B2(new_n260), .ZN(new_n263));
  INV_X1    g062(.A(new_n252), .ZN(new_n264));
  OAI21_X1  g063(.A(G22gat), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G78gat), .B(G106gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT84), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT31), .B(G50gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n262), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n262), .B2(new_n265), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n278), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G127gat), .ZN(new_n286));
  INV_X1    g085(.A(G127gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(KEYINPUT82), .A3(new_n288), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n250), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n210), .A2(new_n214), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n291), .A2(new_n300), .A3(new_n292), .A4(new_n215), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n289), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n301), .A2(new_n303), .A3(new_n297), .A4(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n273), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(G85gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n273), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n315), .B2(new_n306), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n307), .A2(new_n312), .A3(new_n313), .A4(new_n317), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT76), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT66), .B(G183gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(new_n329), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n324), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n333), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(KEYINPUT67), .C1(new_n327), .C2(new_n330), .ZN(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  INV_X1    g137(.A(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT68), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n340), .A2(KEYINPUT26), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(KEYINPUT26), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n341), .B(new_n342), .C1(new_n338), .C2(new_n339), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n334), .A2(new_n335), .A3(new_n337), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT23), .B1(new_n338), .B2(new_n339), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n335), .B(KEYINPUT24), .Z(new_n348));
  NOR2_X1   g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT65), .B(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n351), .A2(new_n352), .A3(G169gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n345), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(G169gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(new_n339), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n326), .A2(G190gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n357), .B(new_n347), .C1(new_n348), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n323), .B1(new_n361), .B2(new_n216), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n322), .B1(new_n344), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n255), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n216), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(new_n322), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n344), .B2(new_n360), .ZN(new_n370));
  INV_X1    g169(.A(new_n322), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT78), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n239), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n361), .A2(new_n323), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n369), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(KEYINPUT77), .B(new_n255), .C1(new_n362), .C2(new_n363), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n380), .B(KEYINPUT79), .Z(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n366), .A2(new_n375), .A3(new_n376), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n384), .A2(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n272), .B1(new_n321), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n361), .A2(new_n289), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n344), .A2(new_n360), .A3(new_n286), .A4(new_n288), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(G227gat), .B2(G233gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT34), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n390), .A2(new_n391), .A3(G227gat), .A4(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G71gat), .B(G99gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT71), .ZN(new_n401));
  XOR2_X1   g200(.A(G15gat), .B(G43gat), .Z(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n395), .B(KEYINPUT32), .C1(new_n398), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n394), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n406), .A3(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT36), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT36), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n393), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n407), .A3(KEYINPUT72), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n307), .A2(new_n312), .A3(new_n313), .A4(new_n317), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n316), .A2(new_n318), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n311), .B(KEYINPUT87), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n315), .A2(new_n306), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n384), .B(new_n420), .C1(new_n421), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n369), .A2(new_n374), .A3(new_n372), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n239), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n255), .A2(new_n362), .A3(new_n363), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(KEYINPUT89), .A3(new_n239), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT37), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n377), .A2(KEYINPUT37), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n381), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n383), .B1(new_n377), .B2(KEYINPUT37), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(KEYINPUT90), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n435), .C1(KEYINPUT90), .C2(new_n439), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n425), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n293), .A2(KEYINPUT88), .A3(new_n297), .A4(new_n295), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n298), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n296), .A2(new_n298), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT39), .B(new_n443), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n449), .A3(new_n298), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n423), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n424), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(KEYINPUT40), .A3(new_n423), .A4(new_n450), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n272), .B1(new_n456), .B2(new_n387), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n389), .B(new_n419), .C1(new_n442), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n420), .B1(new_n421), .B2(new_n424), .ZN(new_n460));
  AND4_X1   g259(.A1(new_n459), .A2(new_n460), .A3(new_n410), .A4(new_n387), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n272), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n415), .A2(new_n416), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n463), .A2(new_n272), .A3(new_n321), .A4(new_n387), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(G29gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT92), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G29gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n472), .A3(G36gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  OR3_X1    g274(.A1(new_n474), .A2(G29gat), .A3(G36gat), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G50gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G43gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G50gat), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT15), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT15), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n477), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n480), .A2(G50gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n478), .A2(G43gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT15), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n476), .A3(new_n475), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT93), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n482), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n498));
  AND2_X1   g297(.A1(G15gat), .A2(G22gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(G15gat), .A2(G22gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G15gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n202), .ZN(new_n503));
  NAND2_X1  g302(.A1(G15gat), .A2(G22gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT94), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507));
  AOI21_X1  g306(.A(G1gat), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT95), .B(new_n509), .C1(new_n501), .C2(new_n505), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n497), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n507), .A3(G1gat), .ZN(new_n517));
  AND4_X1   g316(.A1(new_n497), .A2(new_n516), .A3(new_n517), .A4(new_n513), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n496), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n496), .A2(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n486), .A2(new_n494), .A3(new_n521), .A4(new_n495), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n517), .A3(new_n513), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G8gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n511), .A2(new_n497), .A3(new_n513), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n468), .B(new_n519), .C1(new_n523), .C2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n520), .A2(new_n522), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT96), .A3(new_n468), .A4(new_n519), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n530), .A2(KEYINPUT97), .A3(new_n531), .A4(new_n535), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT11), .B(G169gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT12), .Z(new_n544));
  XOR2_X1   g343(.A(new_n468), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n519), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n527), .A2(new_n496), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n468), .A4(new_n519), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(new_n539), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n550), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n544), .B(KEYINPUT91), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT98), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n551), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n560), .A2(new_n561), .B1(new_n562), .B2(KEYINPUT105), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n562), .B2(KEYINPUT104), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT104), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT105), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT7), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(new_n564), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G99gat), .B(G106gat), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G99gat), .ZN(new_n574));
  INV_X1    g373(.A(G106gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT8), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n566), .A2(new_n571), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n563), .A2(new_n565), .A3(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n578), .B2(new_n570), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G57gat), .B(G64gat), .Z(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  INV_X1    g383(.A(G71gat), .ZN(new_n585));
  INV_X1    g384(.A(G78gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n581), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n579), .A3(new_n590), .A4(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT107), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n594), .A2(new_n593), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(KEYINPUT107), .A3(new_n593), .A4(new_n594), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT108), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n592), .A2(new_n594), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(G230gat), .A3(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT109), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n600), .A2(new_n601), .ZN(new_n613));
  INV_X1    g412(.A(new_n609), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n614), .A3(new_n605), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n559), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n467), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G231gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n242), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT21), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n532), .B1(new_n621), .B2(new_n591), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(G183gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(G183gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n623), .B2(new_n626), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n623), .A2(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n624), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n629), .B1(new_n634), .B2(new_n627), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n620), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n630), .B1(new_n628), .B2(new_n631), .ZN(new_n637));
  INV_X1    g436(.A(new_n620), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n627), .A3(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n591), .A2(new_n621), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT102), .B(G211gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G127gat), .B(G155gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT20), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n644), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n636), .A2(new_n640), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n533), .A2(new_n580), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n653));
  NAND2_X1  g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(new_n496), .ZN(new_n656));
  OAI221_X1 g455(.A(new_n652), .B1(new_n653), .B2(new_n655), .C1(new_n580), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G190gat), .B(G218gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n653), .ZN(new_n663));
  XOR2_X1   g462(.A(G134gat), .B(G162gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n657), .B(new_n658), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT106), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n662), .A2(new_n668), .A3(new_n665), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n618), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n321), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n509), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n387), .ZN(new_n675));
  NAND2_X1  g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n512), .A2(new_n497), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n680), .B(new_n681), .C1(new_n497), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n412), .A2(new_n418), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT110), .B1(new_n411), .B2(new_n417), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n672), .A2(new_n502), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n618), .A2(new_n671), .A3(new_n410), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n502), .B2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n272), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n666), .A2(new_n669), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n458), .B2(new_n466), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n651), .A3(new_n617), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n321), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n470), .A2(new_n472), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n461), .A2(new_n272), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n702));
  INV_X1    g501(.A(new_n425), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT38), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n435), .B1(new_n439), .B2(KEYINPUT90), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n434), .B1(new_n432), .B2(KEYINPUT37), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT38), .B1(new_n708), .B2(new_n381), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n703), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n270), .A2(new_n271), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n712));
  INV_X1    g511(.A(new_n387), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n388), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n702), .B1(new_n715), .B2(new_n686), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n701), .B1(new_n716), .B2(new_n693), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n467), .A2(KEYINPUT44), .A3(new_n670), .ZN(new_n718));
  INV_X1    g517(.A(new_n650), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n647), .B1(new_n636), .B2(new_n640), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n555), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n721), .A2(new_n722), .A3(new_n616), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n717), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n321), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n700), .B1(new_n698), .B2(new_n725), .ZN(G1328gat));
  NOR3_X1   g525(.A1(new_n695), .A2(G36gat), .A3(new_n387), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n724), .B2(new_n387), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1329gat));
  OAI21_X1  g529(.A(G43gat), .B1(new_n724), .B2(new_n686), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n696), .A2(new_n480), .A3(new_n410), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT47), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n711), .A3(new_n718), .A4(new_n723), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n695), .A2(KEYINPUT113), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n272), .A2(G50gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n694), .A2(new_n741), .A3(new_n651), .A4(new_n617), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n738), .A2(new_n743), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(KEYINPUT114), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n744), .A2(KEYINPUT114), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(G1331gat));
  NOR4_X1   g549(.A1(new_n716), .A2(new_n651), .A3(new_n670), .A4(new_n555), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n616), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n697), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756));
  INV_X1    g555(.A(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n713), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT115), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n757), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1333gat));
  INV_X1    g561(.A(new_n410), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n585), .B1(new_n752), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n686), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G71gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n752), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n272), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n586), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n721), .A2(new_n555), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n717), .A2(new_n616), .A3(new_n718), .A4(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n772), .A2(new_n560), .A3(new_n321), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n715), .A2(new_n686), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n670), .B(new_n771), .C1(new_n774), .C2(new_n702), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n697), .A3(new_n616), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n773), .B1(new_n778), .B2(new_n560), .ZN(G1336gat));
  NAND4_X1  g578(.A1(new_n777), .A2(new_n561), .A3(new_n713), .A4(new_n616), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n772), .B2(new_n387), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n781), .B2(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n780), .B(new_n781), .C1(KEYINPUT116), .C2(new_n783), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1337gat));
  NAND4_X1  g586(.A1(new_n777), .A2(new_n574), .A3(new_n410), .A4(new_n616), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n772), .B2(new_n686), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n272), .A2(G106gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n791), .A2(new_n616), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G106gat), .B1(new_n772), .B2(new_n272), .ZN(new_n795));
  NAND2_X1  g594(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n600), .A2(new_n801), .A3(new_n602), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n609), .ZN(new_n803));
  INV_X1    g602(.A(new_n613), .ZN(new_n804));
  INV_X1    g603(.A(new_n602), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n597), .A2(new_n598), .A3(new_n599), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT54), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n613), .A2(new_n809), .A3(KEYINPUT54), .A4(new_n806), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n800), .B(new_n803), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n615), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n810), .ZN(new_n815));
  INV_X1    g614(.A(new_n803), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n814), .B(new_n615), .C1(new_n817), .C2(new_n800), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n800), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n813), .A2(new_n818), .A3(new_n555), .A4(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n543), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n546), .A2(new_n547), .A3(new_n545), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n468), .B1(new_n534), .B2(new_n519), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n551), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n616), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n670), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n813), .A2(new_n818), .A3(new_n825), .A4(new_n819), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n693), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n651), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n616), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n721), .A2(new_n693), .A3(new_n722), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n272), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT120), .A3(new_n272), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(new_n697), .A3(new_n387), .A4(new_n410), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n559), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n321), .B1(new_n830), .B2(new_n832), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n463), .A2(new_n272), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n841), .A2(new_n387), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n276), .A3(new_n555), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n839), .B2(new_n831), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n274), .A3(new_n616), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1341gat));
  XOR2_X1   g648(.A(KEYINPUT69), .B(G127gat), .Z(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n839), .B2(new_n651), .ZN(new_n851));
  INV_X1    g650(.A(new_n844), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(new_n850), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n651), .B2(new_n853), .ZN(G1342gat));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n283), .A3(new_n670), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT56), .Z(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n839), .B2(new_n693), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1343gat));
  NOR2_X1   g657(.A1(new_n765), .A2(new_n272), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT123), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n841), .A2(new_n387), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n559), .A2(G141gat), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT124), .Z(new_n864));
  NOR2_X1   g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n811), .A2(new_n812), .ZN(new_n867));
  XNOR2_X1  g666(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n817), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n556), .A2(new_n558), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n826), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n693), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n828), .A2(new_n693), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n721), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR4_X1   g673(.A1(new_n651), .A2(new_n670), .A3(new_n555), .A4(new_n616), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n711), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n833), .A2(new_n711), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n670), .B1(new_n870), .B2(new_n826), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n651), .B1(new_n882), .B2(new_n829), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(new_n832), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n711), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n878), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n686), .A2(new_n697), .A3(new_n387), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n559), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n866), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n555), .A3(new_n888), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n865), .B1(new_n892), .B2(G141gat), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n879), .A2(KEYINPUT57), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n671), .A2(new_n559), .A3(new_n831), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n880), .B(new_n711), .C1(new_n897), .C2(new_n874), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n616), .A2(new_n896), .A3(new_n898), .A4(new_n888), .ZN(new_n899));
  INV_X1    g698(.A(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n889), .B2(new_n831), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n903), .B2(new_n900), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n860), .A2(new_n900), .A3(new_n861), .A4(new_n616), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1345gat));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n204), .A3(new_n651), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n860), .A2(new_n721), .A3(new_n861), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n204), .B2(new_n908), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n670), .A3(new_n888), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G162gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n860), .A2(new_n205), .A3(new_n861), .A4(new_n670), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n697), .A2(new_n387), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n410), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n836), .A2(new_n837), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n559), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n697), .B1(new_n830), .B2(new_n832), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(new_n713), .A3(new_n843), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n338), .A3(new_n555), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(G1348gat));
  AOI21_X1  g726(.A(G176gat), .B1(new_n925), .B2(new_n616), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n616), .A2(new_n351), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n921), .B2(new_n929), .ZN(G1349gat));
  INV_X1    g729(.A(new_n326), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n921), .B2(new_n721), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n925), .A2(new_n721), .A3(new_n332), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n932), .A2(KEYINPUT60), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT60), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n925), .A2(new_n329), .A3(new_n670), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n836), .A2(new_n670), .A3(new_n837), .A4(new_n920), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G190gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n943), .A3(G190gat), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n941), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(G1351gat));
  NAND4_X1  g746(.A1(new_n896), .A2(new_n898), .A3(new_n686), .A4(new_n918), .ZN(new_n948));
  OAI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n559), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n924), .A2(new_n713), .A3(new_n859), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n219), .A3(new_n555), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(G1352gat));
  OR3_X1    g752(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n831), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n948), .B2(new_n831), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(G204gat), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(new_n220), .A3(new_n616), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  OR3_X1    g759(.A1(new_n950), .A2(G211gat), .A3(new_n651), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n948), .A2(new_n651), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT63), .B(G211gat), .C1(new_n948), .C2(new_n651), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n948), .B2(new_n693), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n950), .A2(G218gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n693), .B2(new_n968), .ZN(G1355gat));
endmodule


