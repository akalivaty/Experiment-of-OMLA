//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT65), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n205), .A2(new_n207), .A3(new_n215), .A4(new_n208), .ZN(new_n216));
  INV_X1    g015(.A(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n211), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n210), .A2(new_n214), .A3(new_n216), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT67), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n212), .A2(new_n213), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n224), .B1(new_n208), .B2(KEYINPUT68), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(new_n230), .A3(new_n207), .A4(new_n205), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n236), .A2(new_n219), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n234), .A2(new_n238), .A3(KEYINPUT28), .A4(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n234), .A2(new_n238), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT28), .A4(new_n219), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT26), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n249), .A2(new_n208), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(KEYINPUT71), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n232), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  INV_X1    g059(.A(new_n254), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT71), .B1(new_n247), .B2(new_n250), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n231), .A2(new_n228), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n223), .A2(new_n224), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n264), .B1(new_n267), .B2(new_n225), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n260), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT77), .A3(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(new_n251), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT78), .B1(new_n272), .B2(new_n257), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(new_n258), .C1(new_n268), .C2(new_n271), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n270), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT76), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(KEYINPUT76), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n277), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288));
  INV_X1    g087(.A(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n257), .B1(new_n272), .B2(KEYINPUT29), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n257), .B1(new_n232), .B2(new_n255), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n291), .A2(KEYINPUT79), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(KEYINPUT79), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n289), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT38), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n276), .A2(new_n289), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n286), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT37), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n276), .A2(new_n289), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT91), .A3(KEYINPUT37), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G141gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT81), .B(G141gat), .Z(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT2), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(KEYINPUT2), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  XNOR2_X1  g120(.A(G155gat), .B(G162gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G155gat), .B(G162gat), .Z(new_n325));
  XNOR2_X1  g124(.A(G141gat), .B(G148gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(KEYINPUT80), .C1(KEYINPUT2), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT2), .B1(new_n312), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G113gat), .B(G120gat), .Z(new_n337));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338));
  INV_X1    g137(.A(G134gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G127gat), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n337), .A2(new_n338), .B1(KEYINPUT72), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g141(.A(G127gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G120gat), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(G113gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT1), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT73), .B1(new_n353), .B2(new_n346), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n345), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n332), .B(new_n327), .C1(new_n315), .C2(new_n323), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT4), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n347), .A2(new_n348), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(KEYINPUT73), .A3(new_n346), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n362), .B1(new_n344), .B2(new_n341), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n334), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n359), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT83), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n310), .B(new_n358), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n355), .B(new_n356), .ZN(new_n370));
  INV_X1    g169(.A(new_n310), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n358), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n364), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n364), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n373), .A2(new_n371), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT86), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n359), .A2(new_n364), .A3(new_n378), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n359), .B2(new_n364), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n358), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n374), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  INV_X1    g188(.A(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT92), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT92), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n388), .A2(new_n396), .A3(KEYINPUT6), .A4(new_n393), .ZN(new_n397));
  INV_X1    g196(.A(new_n393), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n374), .B(new_n398), .C1(new_n382), .C2(new_n387), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT6), .B1(new_n388), .B2(new_n393), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n395), .A2(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n295), .A2(new_n299), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n288), .B1(new_n287), .B2(new_n294), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT38), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n299), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n287), .A2(new_n405), .A3(new_n294), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n309), .A2(new_n401), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  XOR2_X1   g210(.A(new_n411), .B(KEYINPUT89), .Z(new_n412));
  AOI21_X1  g211(.A(new_n289), .B1(new_n336), .B2(new_n260), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G228gat), .ZN(new_n415));
  INV_X1    g214(.A(G233gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n260), .B1(new_n283), .B2(new_n285), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n334), .B1(new_n418), .B2(new_n335), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n413), .A2(new_n419), .B1(new_n415), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G22gat), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n412), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n411), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(KEYINPUT90), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(KEYINPUT90), .A3(G22gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n287), .A2(new_n294), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n299), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n388), .A2(new_n393), .ZN(new_n437));
  OR3_X1    g236(.A1(new_n380), .A2(KEYINPUT39), .A3(new_n310), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n380), .A2(new_n310), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT39), .B1(new_n370), .B2(new_n371), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n438), .B(new_n398), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OR3_X1    g243(.A1(new_n434), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n436), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n407), .A2(new_n433), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n355), .B1(new_n263), .B2(new_n268), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT64), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n232), .A2(new_n255), .A3(new_n363), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT34), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n449), .A2(new_n453), .A3(new_n456), .A4(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(G15gat), .B(G43gat), .Z(new_n460));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n452), .B1(new_n449), .B2(new_n453), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT74), .B(KEYINPUT33), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n453), .ZN(new_n470));
  AOI221_X4 g269(.A(new_n467), .B1(new_n465), .B2(new_n462), .C1(new_n470), .C2(new_n451), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT75), .B(new_n459), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n451), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n464), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n462), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n455), .A2(KEYINPUT75), .A3(new_n457), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n466), .A2(new_n468), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n472), .A2(new_n481), .A3(KEYINPUT36), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n436), .A2(new_n445), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n400), .A2(KEYINPUT87), .A3(new_n399), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n388), .B(new_n393), .C1(new_n489), .C2(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n486), .B1(new_n492), .B2(new_n432), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n432), .B1(new_n472), .B2(new_n481), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  INV_X1    g295(.A(new_n401), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n487), .A3(new_n498), .A4(new_n494), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n448), .A2(new_n493), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G71gat), .ZN(new_n501));
  INV_X1    g300(.A(G78gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT97), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(KEYINPUT97), .A3(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n504), .ZN(new_n510));
  INV_X1    g309(.A(G64gat), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n511), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(G57gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT96), .B1(new_n511), .B2(G57gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n505), .ZN(new_n516));
  XOR2_X1   g315(.A(G57gat), .B(G64gat), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT9), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n510), .A2(new_n515), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT21), .ZN(new_n520));
  XNOR2_X1  g319(.A(G127gat), .B(G155gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G183gat), .B(G211gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT98), .ZN(new_n524));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  XNOR2_X1  g325(.A(new_n522), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT16), .A3(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(new_n529), .C2(new_n528), .ZN(new_n532));
  AND2_X1   g331(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT21), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n510), .A2(new_n515), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n516), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n534), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n527), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT99), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(KEYINPUT41), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT102), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n390), .ZN(new_n555));
  NAND2_X1  g354(.A1(KEYINPUT100), .A2(G85gat), .ZN(new_n556));
  AOI21_X1  g355(.A(G92gat), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT8), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(G99gat), .B2(G106gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  AND2_X1   g360(.A1(KEYINPUT100), .A2(G85gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(KEYINPUT100), .A2(G85gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G99gat), .ZN(new_n565));
  INV_X1    g364(.A(G106gat), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT8), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(KEYINPUT101), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n552), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  AOI211_X1 g373(.A(new_n551), .B(new_n572), .C1(new_n560), .C2(new_n568), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n577));
  INV_X1    g376(.A(G29gat), .ZN(new_n578));
  INV_X1    g377(.A(G36gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n580), .A2(new_n581), .B1(G29gat), .B2(G36gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G43gat), .B(G50gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT15), .ZN(new_n584));
  INV_X1    g383(.A(G43gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(G50gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n586), .B2(KEYINPUT93), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n583), .B1(new_n582), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n547), .A2(KEYINPUT102), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n545), .B2(KEYINPUT41), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n588), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT17), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n597), .A3(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n592), .B(new_n594), .C1(new_n599), .C2(new_n576), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n550), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n549), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n542), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n538), .B1(new_n574), .B2(new_n575), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n564), .A2(KEYINPUT101), .A3(new_n567), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT101), .B1(new_n564), .B2(new_n567), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n573), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n551), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n569), .A2(new_n552), .A3(new_n573), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n519), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n576), .A2(KEYINPUT10), .A3(new_n519), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  AOI211_X1 g423(.A(KEYINPUT105), .B(new_n624), .C1(new_n619), .C2(new_n620), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n617), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT104), .B(G176gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT103), .B1(new_n621), .B2(new_n622), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n637), .B(new_n624), .C1(new_n619), .C2(new_n620), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n628), .B(new_n633), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n596), .A2(new_n534), .A3(new_n598), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n596), .A2(new_n534), .A3(new_n645), .A4(new_n598), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n534), .A2(new_n595), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n643), .A2(new_n644), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n642), .B2(KEYINPUT95), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n652), .A2(KEYINPUT18), .A3(new_n644), .A4(new_n646), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n534), .B(new_n595), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n644), .B(KEYINPUT13), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  INV_X1    g457(.A(G197gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT11), .B(G169gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n651), .A2(new_n653), .A3(new_n656), .A4(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n500), .A2(new_n609), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n491), .B(KEYINPUT106), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  INV_X1    g471(.A(new_n487), .ZN(new_n673));
  NAND2_X1  g472(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n674));
  OR2_X1    g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n669), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n669), .A2(new_n673), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(G8gat), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n676), .B2(new_n680), .ZN(G1325gat));
  AOI21_X1  g480(.A(G15gat), .B1(new_n669), .B2(new_n482), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n486), .A2(G15gat), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n669), .B2(new_n683), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n432), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n448), .A2(new_n493), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n496), .A2(new_n499), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n608), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n668), .A2(new_n542), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n578), .A3(new_n670), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(new_n692), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n500), .B2(new_n608), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  INV_X1    g498(.A(new_n608), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n472), .A2(new_n481), .A3(KEYINPUT36), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT36), .B1(new_n472), .B2(new_n481), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n436), .A2(new_n445), .B1(new_n488), .B2(new_n490), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n433), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n447), .A2(new_n433), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n407), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n487), .A2(new_n494), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n401), .A2(KEYINPUT35), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n709), .A2(new_n710), .B1(new_n495), .B2(KEYINPUT35), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n699), .B(new_n700), .C1(new_n707), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n697), .B1(new_n698), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(new_n670), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n696), .B1(new_n578), .B2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n693), .A2(G36gat), .A3(new_n487), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n713), .A2(new_n718), .A3(new_n673), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G36gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n713), .B2(new_n673), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n694), .A2(new_n585), .A3(new_n482), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n713), .A2(new_n486), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n585), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT47), .B(new_n723), .C1(new_n724), .C2(new_n585), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  AOI211_X1 g528(.A(new_n433), .B(new_n697), .C1(new_n698), .C2(new_n712), .ZN(new_n730));
  INV_X1    g529(.A(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n694), .A2(new_n731), .A3(new_n432), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI221_X1 g535(.A(new_n733), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n730), .C2(new_n731), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n689), .A2(new_n690), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n641), .A2(new_n609), .A3(new_n667), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(KEYINPUT110), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n491), .B(KEYINPUT106), .Z(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(G57gat), .Z(G1332gat));
  OAI22_X1  g547(.A1(new_n745), .A2(new_n487), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n743), .A2(new_n673), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT111), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n755), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n745), .B2(new_n703), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n501), .A3(new_n482), .A4(new_n744), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n433), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n502), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n667), .A2(new_n542), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n691), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n767), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n500), .A2(KEYINPUT51), .A3(new_n608), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n670), .A3(new_n640), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n555), .A2(new_n556), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n641), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n698), .B2(new_n712), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n746), .A2(new_n773), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n772), .A2(new_n773), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  OAI211_X1 g577(.A(new_n700), .B(new_n767), .C1(new_n707), .C2(new_n711), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n768), .B2(new_n770), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(KEYINPUT112), .A3(new_n766), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n487), .A2(G92gat), .A3(new_n641), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n673), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n771), .B2(new_n783), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1337gat));
  NAND3_X1  g590(.A1(new_n771), .A2(new_n482), .A3(new_n640), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n703), .A2(new_n565), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(new_n565), .B1(new_n776), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n433), .A2(G106gat), .A3(new_n641), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n781), .A2(new_n782), .A3(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n433), .B(new_n775), .C1(new_n698), .C2(new_n712), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n566), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT53), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n768), .A2(new_n770), .A3(new_n641), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n433), .A2(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n797), .B2(KEYINPUT113), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n776), .A2(KEYINPUT113), .A3(new_n432), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n805), .ZN(G1339gat));
  INV_X1    g605(.A(new_n542), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n619), .A2(new_n624), .A3(new_n620), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n619), .A2(KEYINPUT114), .A3(new_n620), .A4(new_n624), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(new_n812), .C1(new_n636), .C2(new_n638), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n623), .B2(new_n625), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n634), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT115), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n814), .A4(new_n634), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n639), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(new_n821), .A3(new_n816), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n818), .A2(new_n820), .A3(new_n667), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n644), .B1(new_n652), .B2(new_n646), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n654), .A2(new_n655), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n662), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n666), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n640), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n700), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n822), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n821), .B1(new_n815), .B2(new_n816), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n819), .A2(new_n639), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n607), .A2(new_n605), .A3(new_n666), .A4(new_n826), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n807), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n609), .A2(new_n640), .A3(new_n667), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n670), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n708), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n667), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g641(.A(new_n350), .B1(new_n840), .B2(new_n640), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT116), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n640), .A2(new_n350), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT117), .Z(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(G1341gat));
  NAND2_X1  g647(.A1(new_n840), .A2(new_n542), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n840), .A2(new_n700), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n339), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n339), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(KEYINPUT56), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(KEYINPUT56), .B2(new_n854), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n746), .B1(new_n835), .B2(new_n837), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n486), .A2(new_n433), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n673), .B1(new_n862), .B2(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n667), .A2(new_n329), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n858), .A2(new_n866), .A3(new_n860), .A4(new_n861), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n861), .B1(new_n859), .B2(KEYINPUT118), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n838), .A2(KEYINPUT118), .A3(new_n670), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n867), .A3(new_n487), .A4(new_n865), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n433), .B1(new_n835), .B2(new_n837), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n815), .A2(new_n816), .B1(new_n665), .B2(new_n666), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n820), .A2(new_n878), .B1(new_n640), .B2(new_n827), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n818), .A2(new_n820), .A3(new_n822), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n879), .A2(new_n700), .B1(new_n880), .B2(new_n833), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n836), .B1(new_n881), .B2(new_n807), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n433), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n746), .A2(new_n673), .A3(new_n486), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n877), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n314), .B1(new_n885), .B2(new_n667), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT58), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n874), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n862), .A2(new_n673), .A3(new_n864), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n432), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n817), .A2(new_n667), .A3(new_n639), .A4(new_n819), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n700), .B1(new_n894), .B2(new_n828), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n807), .B1(new_n834), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n433), .B1(new_n896), .B2(new_n837), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT121), .B1(new_n897), .B2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n899), .B(new_n876), .C1(new_n882), .C2(new_n433), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n640), .A3(new_n884), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n311), .B1(new_n902), .B2(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n901), .A2(new_n904), .A3(new_n640), .A4(new_n884), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n892), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n311), .C1(new_n885), .C2(new_n640), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n863), .A2(new_n867), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n640), .A2(new_n311), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1345gat));
  NAND3_X1  g709(.A1(new_n863), .A2(new_n542), .A3(new_n867), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n807), .A2(new_n316), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n911), .A2(new_n316), .B1(new_n885), .B2(new_n912), .ZN(G1346gat));
  NAND2_X1  g712(.A1(new_n700), .A2(new_n317), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n885), .A2(new_n700), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n908), .A2(new_n914), .B1(new_n317), .B2(new_n915), .ZN(G1347gat));
  NAND2_X1  g715(.A1(new_n673), .A2(new_n494), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n670), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n838), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n667), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(G169gat), .ZN(G1348gat));
  NOR2_X1   g721(.A1(new_n919), .A2(new_n641), .ZN(new_n923));
  XOR2_X1   g722(.A(KEYINPUT123), .B(G176gat), .Z(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n920), .A2(new_n542), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n218), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n926), .B2(new_n244), .ZN(new_n928));
  XNOR2_X1  g727(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1350gat));
  NOR2_X1   g729(.A1(new_n919), .A2(new_n608), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n219), .ZN(new_n933));
  XOR2_X1   g732(.A(KEYINPUT61), .B(G190gat), .Z(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n931), .B2(new_n934), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n670), .A2(new_n487), .A3(new_n486), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n875), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n659), .A3(new_n667), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n901), .A2(new_n667), .A3(new_n936), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G197gat), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  INV_X1    g742(.A(G204gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n937), .A2(new_n944), .A3(new_n640), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT62), .Z(new_n946));
  AND3_X1   g745(.A1(new_n901), .A2(new_n640), .A3(new_n936), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n944), .B2(new_n947), .ZN(G1353gat));
  INV_X1    g747(.A(G211gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n949), .A3(new_n542), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n901), .A2(new_n542), .A3(new_n936), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G211gat), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(KEYINPUT126), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT126), .B1(new_n952), .B2(new_n953), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n950), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n937), .A2(new_n959), .A3(new_n700), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n901), .A2(KEYINPUT127), .A3(new_n936), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT127), .B1(new_n901), .B2(new_n936), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n608), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n963), .B2(new_n959), .ZN(G1355gat));
endmodule


