//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(G355));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  AND2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT67), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n204), .A2(new_n205), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n223), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G58), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI211_X1 g0054(.A(G1), .B(G13), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n253), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G226), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT72), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT72), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n262), .A3(G226), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n257), .A2(new_n258), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G232), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n255), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n255), .A2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(G238), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT13), .B1(new_n271), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n269), .B1(new_n263), .B2(new_n261), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n279), .C1(new_n283), .C2(new_n255), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G190), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT73), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT73), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n281), .A2(new_n287), .A3(G190), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n230), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n274), .A2(G20), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n294), .A2(G68), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n231), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n228), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(new_n293), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n296), .B1(new_n303), .B2(KEYINPUT11), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT74), .B1(new_n290), .B2(G68), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n305), .B(KEYINPUT12), .Z(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n306), .C1(KEYINPUT11), .C2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n281), .A2(new_n284), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(G200), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n289), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n281), .A2(G179), .A3(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n281), .A2(KEYINPUT75), .A3(G179), .A4(new_n284), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n308), .A2(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(new_n318), .A3(G169), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n307), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n274), .B2(G20), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n294), .A2(new_n324), .B1(new_n323), .B2(new_n291), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n298), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n300), .B1(G20), .B2(G77), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n326), .B1(new_n338), .B2(new_n293), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n292), .A2(new_n230), .ZN(new_n340));
  AOI211_X1 g0140(.A(KEYINPUT70), .B(new_n340), .C1(new_n332), .C2(new_n337), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n325), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n275), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n255), .A3(G274), .ZN(new_n344));
  INV_X1    g0144(.A(G244), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n277), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G107), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n347), .B(new_n351), .C1(new_n267), .C2(G1698), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n272), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(G169), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n342), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(G190), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n353), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n342), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n322), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n259), .A2(G222), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n266), .A2(G223), .A3(G1698), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n364), .C1(new_n323), .C2(new_n266), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n272), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n344), .B1(new_n277), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(G179), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n231), .B1(new_n227), .B2(new_n228), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT8), .B(G58), .ZN(new_n373));
  INV_X1    g0173(.A(G150), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n297), .B1(new_n374), .B2(new_n301), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n293), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n228), .B1(new_n274), .B2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n294), .A2(new_n377), .B1(new_n228), .B2(new_n291), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n368), .B1(new_n365), .B2(new_n272), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(G169), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n371), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n370), .A2(new_n384), .B1(new_n380), .B2(KEYINPUT9), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT9), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n381), .A2(new_n359), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT10), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT10), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n381), .A2(G190), .B1(new_n379), .B2(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n383), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n342), .A2(new_n360), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n342), .A2(new_n354), .A3(new_n356), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n362), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n257), .A2(new_n231), .A3(new_n258), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n258), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(G68), .ZN(new_n406));
  AOI211_X1 g0206(.A(KEYINPUT76), .B(new_n203), .C1(new_n403), .C2(new_n404), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n399), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n350), .B2(new_n231), .ZN(new_n409));
  INV_X1    g0209(.A(new_n404), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n399), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n340), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n367), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n266), .B(new_n417), .C1(G223), .C2(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n255), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n344), .B1(new_n277), .B2(new_n237), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n359), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n418), .A2(new_n419), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n255), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(G190), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n340), .A2(new_n290), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n336), .A2(new_n295), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n290), .B2(new_n336), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT77), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n415), .A2(new_n416), .A3(new_n426), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n415), .A2(new_n432), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n420), .A2(new_n355), .A3(new_n421), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n425), .B2(G169), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n431), .B1(new_n408), .B2(new_n414), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(new_n416), .A3(KEYINPUT17), .A4(new_n426), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT18), .B1(new_n442), .B2(new_n439), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n435), .A2(new_n441), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n310), .A2(new_n321), .A3(new_n397), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n266), .A2(G264), .A3(G1698), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n266), .A2(G257), .A3(new_n268), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT81), .B(G303), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n350), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n272), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G1), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n272), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n455), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n272), .A2(new_n273), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n457), .A2(G270), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n274), .A2(G33), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n294), .A2(G116), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n292), .A2(new_n230), .B1(G20), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n231), .C1(G33), .C2(new_n207), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT20), .B1(new_n465), .B2(new_n467), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n463), .B1(G116), .B2(new_n290), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n461), .A2(new_n470), .A3(G169), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n461), .A2(new_n355), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n472), .A2(KEYINPUT21), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(KEYINPUT82), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n470), .B1(new_n461), .B2(G200), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n384), .B2(new_n461), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n474), .A2(new_n481), .A3(new_n476), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n484));
  OAI211_X1 g0284(.A(G244), .B(new_n268), .C1(new_n348), .C2(new_n349), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n466), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT4), .B1(new_n259), .B2(G244), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n272), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n457), .A2(G257), .B1(new_n458), .B2(new_n459), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT79), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(KEYINPUT79), .A3(new_n490), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(G190), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT6), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n496), .A2(new_n207), .A3(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(G97), .B(G107), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n499), .A2(new_n231), .B1(new_n323), .B2(new_n301), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n208), .B1(new_n403), .B2(new_n404), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n293), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n290), .A2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n294), .A2(new_n462), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n491), .A2(G200), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n495), .A2(new_n502), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n456), .A2(new_n455), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(G264), .A3(new_n255), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT85), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n457), .A2(new_n512), .A3(G264), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n458), .A2(new_n459), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n259), .A2(G250), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n259), .A2(KEYINPUT84), .A3(G250), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n514), .B(new_n515), .C1(new_n523), .C2(new_n255), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n516), .A2(new_n517), .ZN(new_n526));
  INV_X1    g0326(.A(new_n522), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT84), .B1(new_n259), .B2(G250), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n272), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(G190), .A3(new_n515), .A4(new_n514), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n266), .A2(new_n231), .A3(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n266), .A2(new_n534), .A3(new_n231), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n231), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n537), .B1(new_n536), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n293), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT25), .B1(new_n291), .B2(new_n208), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n505), .A2(G107), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n525), .A2(new_n531), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n266), .A2(G244), .A3(G1698), .ZN(new_n552));
  OAI211_X1 g0352(.A(G238), .B(new_n268), .C1(new_n348), .C2(new_n349), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n538), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n272), .ZN(new_n555));
  OR3_X1    g0355(.A1(new_n454), .A2(KEYINPUT80), .A3(G1), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT80), .B1(new_n454), .B2(G1), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n255), .A2(G250), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n459), .B2(new_n455), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n266), .A2(new_n231), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n231), .B1(new_n265), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G87), .B2(new_n209), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n297), .B2(new_n207), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n293), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n328), .A2(new_n331), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n291), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n294), .A2(G87), .A3(new_n462), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n555), .A2(new_n560), .A3(G190), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n562), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n328), .A2(new_n294), .A3(new_n331), .A4(new_n462), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n555), .A2(new_n560), .A3(new_n355), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n459), .A2(new_n455), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n556), .A2(new_n255), .A3(new_n557), .A4(G250), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n272), .B2(new_n554), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n577), .B(new_n578), .C1(new_n582), .C2(G169), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G169), .ZN(new_n585));
  INV_X1    g0385(.A(new_n494), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT79), .B1(new_n489), .B2(new_n490), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n491), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n355), .B1(new_n502), .B2(new_n506), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n508), .A2(new_n551), .A3(new_n584), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n524), .A2(new_n585), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n530), .A2(new_n355), .A3(new_n515), .A4(new_n514), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n536), .A2(new_n543), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n340), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n550), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n447), .A2(new_n483), .A3(new_n602), .ZN(G372));
  NAND4_X1  g0403(.A1(new_n588), .A2(new_n590), .A3(new_n583), .A4(new_n575), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT26), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n474), .A2(new_n600), .A3(new_n476), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n583), .B1(new_n606), .B2(new_n592), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n447), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n383), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n441), .A2(new_n444), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n289), .A2(new_n309), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n321), .B1(new_n611), .B2(new_n395), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n435), .A2(new_n443), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n388), .A2(new_n392), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(KEYINPUT86), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n608), .B(new_n609), .C1(new_n615), .C2(new_n619), .ZN(G369));
  AND2_X1   g0420(.A1(new_n480), .A2(new_n482), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT88), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n274), .A2(new_n231), .A3(G13), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n470), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT87), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n483), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n474), .A2(new_n476), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n600), .A2(new_n628), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n628), .B1(new_n598), .B2(new_n599), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n551), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n637), .B1(new_n600), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(G330), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n635), .A2(new_n628), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n600), .B2(new_n628), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(G399));
  INV_X1    g0446(.A(new_n224), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G41), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G1), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n229), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT31), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n514), .B1(new_n523), .B2(new_n255), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT89), .B1(new_n656), .B2(new_n561), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n530), .A2(new_n582), .A3(new_n658), .A4(new_n514), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n473), .A2(new_n493), .A3(new_n494), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(KEYINPUT30), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(G179), .B1(new_n453), .B2(new_n460), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n524), .A2(new_n664), .A3(new_n491), .A4(new_n561), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT30), .B1(new_n660), .B2(new_n661), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n628), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n655), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n483), .A2(new_n602), .A3(new_n668), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n666), .A2(new_n665), .ZN(new_n671));
  OAI211_X1 g0471(.A(KEYINPUT31), .B(new_n628), .C1(new_n671), .C2(new_n663), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n668), .B1(new_n607), .B2(new_n605), .ZN(new_n678));
  AND2_X1   g0478(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n682));
  OAI221_X1 g0482(.A(new_n668), .B1(new_n682), .B2(new_n679), .C1(new_n607), .C2(new_n605), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n654), .B1(new_n686), .B2(G1), .ZN(G364));
  NOR2_X1   g0487(.A1(new_n231), .A2(G179), .ZN(new_n688));
  NOR2_X1   g0488(.A1(G190), .A2(G200), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G159), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT32), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n231), .A2(new_n355), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT92), .Z(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(G190), .A3(G200), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n350), .B(new_n693), .C1(new_n696), .C2(G77), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n384), .A3(G200), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n202), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n355), .A2(new_n359), .A3(G190), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G20), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n207), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n694), .A2(G200), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(G68), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n705), .A2(new_n384), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n688), .A2(new_n384), .A3(G200), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n710), .A2(G50), .B1(new_n712), .B2(G107), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n688), .A2(G190), .A3(G200), .ZN(new_n714));
  INV_X1    g0514(.A(G87), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n692), .B2(KEYINPUT32), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n708), .A2(new_n709), .A3(new_n713), .A4(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n710), .A2(G326), .B1(new_n702), .B2(G294), .ZN(new_n719));
  INV_X1    g0519(.A(G317), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT33), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n720), .A2(KEYINPUT33), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n706), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G283), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n719), .B(new_n723), .C1(new_n724), .C2(new_n711), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n266), .B1(new_n691), .B2(G329), .ZN(new_n726));
  INV_X1    g0526(.A(G303), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n714), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n698), .B2(G322), .ZN(new_n729));
  INV_X1    g0529(.A(G311), .ZN(new_n730));
  INV_X1    g0530(.A(new_n696), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n700), .A2(new_n718), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n230), .B1(G20), .B2(new_n585), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n231), .A2(G13), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n274), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n648), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT91), .Z(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n734), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n224), .A2(G355), .A3(new_n266), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n647), .A2(new_n266), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G45), .B2(new_n652), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n251), .A2(new_n454), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n746), .B1(G116), .B2(new_n224), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n741), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n744), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n735), .B(new_n751), .C1(new_n636), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n739), .ZN(new_n754));
  INV_X1    g0554(.A(new_n636), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(new_n675), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n636), .A2(G330), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(G396));
  NOR2_X1   g0558(.A1(new_n734), .A2(new_n742), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n740), .B1(G77), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n706), .ZN(new_n762));
  INV_X1    g0562(.A(new_n710), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n724), .B1(new_n763), .B2(new_n727), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n715), .A2(new_n711), .B1(new_n714), .B2(new_n208), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n266), .B(new_n704), .C1(G311), .C2(new_n691), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n698), .A2(G294), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n696), .A2(G116), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G137), .A2(new_n710), .B1(new_n706), .B2(G150), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  INV_X1    g0572(.A(G143), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n771), .B1(new_n731), .B2(new_n772), .C1(new_n773), .C2(new_n699), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT34), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G132), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n266), .B1(new_n690), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n712), .A2(G68), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n228), .B2(new_n714), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G58), .C2(new_n702), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n774), .A2(new_n775), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n770), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n761), .B1(new_n784), .B2(new_n734), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n395), .A2(new_n628), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n342), .A2(new_n628), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n394), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n395), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n785), .B1(new_n789), .B2(new_n743), .ZN(new_n790));
  INV_X1    g0590(.A(new_n678), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n789), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n668), .B(new_n789), .C1(new_n607), .C2(new_n605), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n792), .B(new_n794), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n754), .B1(new_n796), .B2(new_n676), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n677), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(G384));
  INV_X1    g0599(.A(new_n499), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT35), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(KEYINPUT35), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n801), .A2(G116), .A3(new_n232), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT36), .Z(new_n804));
  OAI211_X1 g0604(.A(new_n229), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n228), .A2(G68), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n274), .B(G13), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT39), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT37), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n442), .A2(new_n426), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n429), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n399), .B1(new_n406), .B2(new_n407), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n340), .B1(new_n814), .B2(new_n413), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n408), .B1(new_n815), .B2(KEYINPUT97), .ZN(new_n816));
  INV_X1    g0616(.A(new_n399), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n411), .A2(KEYINPUT76), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n405), .A2(new_n400), .A3(G68), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(KEYINPUT97), .B(new_n293), .C1(new_n820), .C2(KEYINPUT16), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n813), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n626), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n812), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n440), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n810), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n812), .B1(new_n436), .B2(new_n440), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n436), .A2(KEYINPUT99), .A3(new_n824), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT99), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n442), .B2(new_n626), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n828), .A2(new_n832), .A3(new_n810), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n293), .B1(new_n820), .B2(KEYINPUT16), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT97), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n408), .A3(new_n821), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n626), .B1(new_n837), .B2(new_n813), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT98), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n838), .A2(new_n445), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n838), .B2(new_n445), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n827), .A2(new_n833), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n834), .A2(new_n835), .B1(KEYINPUT16), .B2(new_n820), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n429), .B1(new_n845), .B2(new_n821), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n811), .B1(new_n846), .B2(new_n626), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n439), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n828), .A2(new_n832), .A3(new_n810), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n841), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n838), .A2(new_n445), .A3(new_n839), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n854), .A3(KEYINPUT38), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n844), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n842), .A2(KEYINPUT100), .A3(new_n843), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n809), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n842), .A2(new_n843), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n828), .A2(new_n832), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n850), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n445), .A2(new_n831), .A3(new_n829), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n320), .A2(new_n307), .A3(new_n668), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT101), .Z(new_n869));
  NOR3_X1   g0669(.A1(new_n859), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n610), .A2(new_n626), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n786), .B(KEYINPUT95), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n307), .A2(new_n628), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n321), .A2(new_n310), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n307), .B(new_n628), .C1(new_n611), .C2(new_n320), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n793), .A2(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT96), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n857), .A2(new_n858), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n609), .B1(new_n615), .B2(new_n619), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n681), .A2(new_n447), .A3(new_n683), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n681), .A2(new_n447), .A3(new_n683), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n880), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n874), .A2(new_n875), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n673), .A2(new_n789), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT40), .B1(new_n866), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(KEYINPUT40), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n858), .A3(new_n857), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n673), .A2(new_n447), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n675), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n887), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n274), .B2(new_n736), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n887), .A2(new_n896), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n808), .B1(new_n898), .B2(new_n899), .ZN(G367));
  INV_X1    g0700(.A(new_n747), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n745), .B1(new_n224), .B2(new_n570), .C1(new_n901), .C2(new_n243), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n740), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n573), .A2(new_n668), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT103), .Z(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n584), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n583), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n702), .A2(G68), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n699), .B2(new_n374), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT109), .Z(new_n911));
  INV_X1    g0711(.A(G137), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n266), .B1(new_n690), .B2(new_n912), .C1(new_n762), .C2(new_n772), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n696), .B2(G50), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n711), .A2(new_n323), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G143), .B2(new_n710), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n916), .C1(new_n202), .C2(new_n714), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n350), .B1(new_n690), .B2(new_n720), .C1(new_n207), .C2(new_n711), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n698), .B2(new_n450), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n724), .B2(new_n731), .ZN(new_n920));
  INV_X1    g0720(.A(new_n714), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G116), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n706), .A2(G294), .B1(new_n702), .B2(G107), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n730), .C2(new_n763), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n911), .A2(new_n917), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT47), .Z(new_n927));
  INV_X1    g0727(.A(new_n734), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n903), .B1(new_n752), .B2(new_n908), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n737), .B(KEYINPUT108), .Z(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT107), .B1(new_n640), .B2(new_n642), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n755), .B2(new_n675), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n636), .A2(G330), .A3(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n643), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n643), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n686), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n591), .A2(new_n668), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n508), .A2(new_n591), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n502), .A2(new_n506), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n628), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n644), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT45), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n644), .A2(new_n946), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT44), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n636), .A2(KEYINPUT106), .A3(G330), .A4(new_n640), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n686), .B1(new_n940), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n648), .B(new_n955), .Z(new_n956));
  AOI21_X1  g0756(.A(new_n930), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n643), .A2(new_n946), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n601), .A2(new_n508), .B1(new_n588), .B2(new_n590), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n628), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n908), .B(KEYINPUT43), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n961), .A2(KEYINPUT43), .A3(new_n908), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT104), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n641), .A2(new_n946), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(new_n969), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n929), .B1(new_n957), .B2(new_n970), .ZN(G387));
  OR3_X1    g0771(.A1(new_n240), .A2(new_n454), .A3(new_n266), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n373), .A2(G50), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n974));
  OAI221_X1 g0774(.A(new_n454), .B1(new_n203), .B2(new_n323), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n350), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n650), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n647), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n745), .B1(new_n224), .B2(new_n208), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n740), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT112), .Z(new_n982));
  AOI22_X1  g0782(.A1(new_n696), .A2(G68), .B1(new_n336), .B2(new_n706), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT113), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n266), .B1(new_n690), .B2(new_n374), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n763), .A2(new_n772), .B1(new_n714), .B2(new_n323), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G97), .C2(new_n712), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n698), .A2(G50), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n328), .A2(new_n331), .A3(new_n702), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n984), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G317), .A2(new_n698), .B1(new_n696), .B2(new_n450), .ZN(new_n991));
  INV_X1    g0791(.A(G322), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n762), .A2(new_n730), .B1(new_n763), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT114), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT48), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(G294), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n703), .A2(new_n724), .B1(new_n714), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n266), .B1(new_n691), .B2(G326), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n464), .B2(new_n711), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT49), .B1(new_n998), .B2(new_n1001), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n990), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n982), .B1(new_n1008), .B2(new_n734), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n640), .B2(new_n752), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT116), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT110), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n939), .B2(new_n930), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n930), .ZN(new_n1014));
  AOI211_X1 g0814(.A(KEYINPUT110), .B(new_n1014), .C1(new_n937), .C2(new_n938), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n648), .B(KEYINPUT117), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n940), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n939), .A2(new_n686), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1011), .B1(new_n1013), .B2(new_n1015), .C1(new_n1017), .C2(new_n1018), .ZN(G393));
  NAND2_X1  g0819(.A1(new_n248), .A2(new_n747), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n745), .C1(new_n207), .C2(new_n224), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n350), .B1(new_n690), .B2(new_n992), .C1(new_n208), .C2(new_n711), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n706), .A2(new_n450), .B1(new_n702), .B2(G116), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n731), .B2(new_n999), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT119), .Z(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(G283), .C2(new_n921), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n698), .A2(G311), .B1(G317), .B2(new_n710), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT52), .Z(new_n1028));
  AOI22_X1  g0828(.A1(new_n698), .A2(G159), .B1(G150), .B2(new_n710), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT51), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n266), .B1(new_n690), .B2(new_n773), .C1(new_n715), .C2(new_n711), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n702), .A2(G77), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n203), .B2(new_n714), .C1(new_n762), .C2(new_n228), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(new_n336), .C2(new_n696), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1026), .A2(new_n1028), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n740), .B(new_n1021), .C1(new_n1035), .C2(new_n928), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n946), .B2(new_n744), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n951), .A2(new_n641), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n951), .A2(new_n641), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT118), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1014), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT118), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n940), .A2(new_n1040), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1016), .B1(new_n940), .B2(new_n953), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G390));
  NAND2_X1  g0847(.A1(new_n676), .A2(new_n447), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n886), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT122), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n886), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n673), .A2(G330), .A3(new_n789), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n888), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n673), .A2(G330), .A3(new_n888), .A4(new_n789), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n793), .A2(new_n872), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n793), .A3(new_n872), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1050), .A2(new_n1052), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1056), .A2(KEYINPUT121), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1056), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT121), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1058), .A2(new_n888), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT120), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n869), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n868), .B(KEYINPUT101), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT120), .B1(new_n876), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n856), .B1(new_n842), .B2(new_n843), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT38), .B1(new_n851), .B2(new_n854), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n858), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT39), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n860), .A2(new_n865), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n809), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1074), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n866), .A2(new_n1072), .A3(new_n876), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1064), .B(new_n1068), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n859), .B2(new_n867), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1083), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1086), .A2(new_n1066), .A3(new_n1065), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1062), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1016), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1062), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n930), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n742), .B1(new_n859), .B2(new_n867), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n741), .B1(new_n373), .B2(new_n759), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n350), .B1(new_n690), .B2(new_n999), .C1(new_n715), .C2(new_n714), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n779), .B1(new_n763), .B2(new_n724), .C1(new_n208), .C2(new_n762), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G97), .C2(new_n696), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1032), .B1(new_n699), .B2(new_n464), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT124), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n350), .B1(new_n691), .B2(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n228), .B2(new_n711), .C1(new_n699), .C2(new_n777), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT123), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n696), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n710), .A2(G128), .B1(new_n702), .B2(G159), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n912), .B2(new_n762), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n714), .B2(new_n374), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n921), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1100), .A2(new_n1102), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1096), .B(new_n1097), .C1(new_n928), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1094), .A2(new_n1095), .A3(new_n1115), .ZN(G378));
  OAI22_X1  g0916(.A1(new_n762), .A2(new_n777), .B1(new_n703), .B2(new_n374), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n698), .A2(G128), .B1(new_n921), .B2(new_n1106), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n696), .A2(G137), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1117), .B(new_n1120), .C1(G125), .C2(new_n710), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n712), .A2(G159), .ZN(new_n1124));
  AOI211_X1 g0924(.A(G33), .B(G41), .C1(new_n691), .C2(G124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT59), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n1121), .ZN(new_n1128));
  AOI211_X1 g0928(.A(G41), .B(new_n266), .C1(new_n691), .C2(G283), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(new_n909), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n731), .B2(new_n570), .C1(new_n208), .C2(new_n699), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n762), .A2(new_n207), .B1(new_n323), .B2(new_n714), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n763), .A2(new_n464), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n711), .A2(new_n202), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT58), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT58), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n266), .A2(G41), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n734), .B1(new_n1128), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n739), .C1(G50), .C2(new_n760), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n617), .A2(new_n609), .A3(new_n618), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n380), .A2(new_n626), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n1151), .B2(new_n742), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n893), .B2(G330), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n893), .A2(new_n1153), .A3(G330), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n880), .A3(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n675), .B(new_n1151), .C1(new_n892), .C2(new_n890), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1158), .A2(new_n1154), .B1(new_n870), .B2(new_n879), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1152), .B1(new_n1160), .B2(new_n930), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1063), .B(new_n1067), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1163));
  AND4_X1   g0963(.A1(new_n1066), .A2(new_n1086), .A3(new_n1065), .A4(new_n1087), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1093), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1168), .B2(KEYINPUT125), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT125), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT125), .B1(new_n1089), .B2(new_n1166), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1171), .A2(new_n1173), .A3(KEYINPUT57), .A4(new_n1160), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1016), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1161), .B1(new_n1172), .B2(new_n1175), .ZN(G375));
  INV_X1    g0976(.A(new_n1061), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n956), .A3(new_n1062), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1061), .A2(new_n930), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n740), .B1(G68), .B2(new_n760), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G107), .A2(new_n696), .B1(new_n698), .B2(G283), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n762), .A2(new_n464), .B1(new_n763), .B2(new_n999), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G97), .B2(new_n921), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n266), .B(new_n915), .C1(G303), .C2(new_n691), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n989), .A4(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n696), .A2(G150), .B1(new_n706), .B2(new_n1106), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n350), .B(new_n1134), .C1(G128), .C2(new_n691), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n912), .C2(new_n699), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n710), .A2(G132), .B1(new_n702), .B2(G50), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n772), .B2(new_n714), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1181), .B1(new_n734), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n888), .B2(new_n743), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1180), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1179), .A2(new_n1196), .ZN(G381));
  OR3_X1    g0997(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1198));
  OR2_X1    g0998(.A1(G393), .A2(G396), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(G387), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(G378), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1161), .A4(new_n1202), .ZN(G407));
  NAND2_X1  g1003(.A1(new_n627), .A2(G213), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G407), .B(G213), .C1(G375), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT126), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1207), .B(new_n1208), .ZN(G409));
  NAND2_X1  g1009(.A1(new_n1205), .A2(G2897), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1178), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n1177), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1016), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT127), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1090), .B1(new_n1212), .B2(new_n1178), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT127), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1214), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1195), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G384), .ZN(new_n1221));
  INV_X1    g1021(.A(G384), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1222), .B(new_n1195), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1211), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1219), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1218), .B1(new_n1217), .B2(new_n1214), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1196), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1222), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1220), .A2(G384), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1210), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1161), .C1(new_n1172), .C2(new_n1175), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1171), .A2(new_n1173), .A3(new_n1160), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n956), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1161), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1201), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1204), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G387), .B(G390), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(G396), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1205), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1242), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1240), .A2(new_n1244), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1248), .A2(new_n1251), .A3(new_n1242), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1248), .B2(new_n1231), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1251), .B1(new_n1248), .B2(new_n1242), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1250), .B1(new_n1256), .B2(new_n1247), .ZN(G405));
  INV_X1    g1057(.A(new_n1247), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(new_n1201), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1233), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1242), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1243), .A3(new_n1233), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1258), .B(new_n1263), .ZN(G402));
endmodule


