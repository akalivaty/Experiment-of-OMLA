//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT77), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n191), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT76), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n190), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  AOI211_X1 g013(.A(KEYINPUT77), .B(new_n199), .C1(new_n194), .C2(new_n196), .ZN(new_n200));
  OAI21_X1  g014(.A(G146), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G237), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G214), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n204), .B(G143), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT90), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT19), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n194), .A2(new_n196), .B1(new_n212), .B2(KEYINPUT90), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(new_n214), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n201), .B(new_n211), .C1(new_n217), .C2(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n208), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n206), .A2(KEYINPUT18), .A3(G131), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n197), .B2(new_n222), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n229), .B(KEYINPUT91), .ZN(new_n232));
  INV_X1    g046(.A(new_n190), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n188), .A2(KEYINPUT76), .A3(G125), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n212), .B2(new_n193), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n235), .B2(new_n199), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT77), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n197), .A2(new_n237), .A3(KEYINPUT16), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n222), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n201), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n207), .A2(new_n210), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n245), .B2(KEYINPUT92), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n225), .B(new_n232), .C1(new_n242), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  NOR2_X1   g063(.A1(G475), .A2(G902), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT93), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n248), .A2(new_n253), .A3(new_n249), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n250), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT20), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G122), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G116), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT14), .ZN(new_n261));
  OR3_X1    g075(.A1(new_n258), .A2(KEYINPUT14), .A3(G116), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(G116), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT94), .A4(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(G107), .C1(KEYINPUT94), .C2(new_n262), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n260), .A2(new_n263), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n205), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n205), .A2(G128), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n265), .B(new_n268), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n266), .B(new_n267), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n277), .B(KEYINPUT13), .Z(new_n283));
  OAI21_X1  g097(.A(G134), .B1(new_n283), .B2(new_n274), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  INV_X1    g101(.A(G217), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n287), .A2(new_n288), .A3(G953), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(new_n285), .A3(new_n289), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G478), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT15), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(KEYINPUT15), .B2(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(G234), .A2(G237), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(G952), .A3(new_n203), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(G902), .A3(G953), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n298), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n225), .B1(new_n242), .B2(new_n246), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n230), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n247), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n294), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G475), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n257), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G221), .B1(new_n287), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT84), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n267), .A3(G104), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n228), .A2(G107), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n228), .A2(G107), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n267), .A2(G104), .ZN(new_n326));
  OAI21_X1  g140(.A(G101), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n222), .A2(G143), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n205), .A2(G146), .ZN(new_n330));
  AND4_X1   g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(G128), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(G128), .B1(new_n329), .B2(new_n330), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n324), .B(new_n327), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n205), .A2(KEYINPUT64), .A3(G146), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n329), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT65), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT0), .A2(G128), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT0), .A2(G128), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n205), .A2(G146), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n222), .B2(G143), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n205), .A2(KEYINPUT64), .A3(G146), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n343), .A2(new_n344), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT65), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n329), .A2(new_n330), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT66), .A3(new_n343), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n329), .A2(new_n330), .A3(new_n343), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n364), .A3(G101), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n354), .A2(new_n357), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n349), .A2(new_n350), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n368), .A2(new_n329), .B1(new_n273), .B2(new_n332), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n369), .B2(new_n331), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n328), .A3(G128), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n273), .A2(new_n332), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(KEYINPUT69), .C1(new_n372), .C2(new_n351), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n324), .A2(new_n327), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n335), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n334), .A2(KEYINPUT82), .A3(new_n335), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n338), .A2(new_n366), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n276), .B2(G137), .ZN(new_n380));
  INV_X1    g194(.A(G137), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT11), .A3(G134), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n276), .A2(G137), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G131), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n382), .A3(new_n209), .A4(new_n383), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G140), .ZN(new_n392));
  INV_X1    g206(.A(G227), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n390), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n371), .B1(new_n372), .B2(new_n351), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n324), .A2(new_n327), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n334), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n400), .A2(KEYINPUT12), .A3(new_n390), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT12), .B1(new_n400), .B2(new_n390), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n378), .A2(new_n390), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n395), .B(KEYINPUT81), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n396), .A2(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT83), .B(G469), .C1(new_n405), .C2(G902), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n407));
  NAND2_X1  g221(.A1(G469), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n334), .A2(KEYINPUT82), .A3(new_n335), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT82), .B1(new_n334), .B2(new_n335), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n390), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n366), .A4(new_n376), .ZN(new_n414));
  INV_X1    g228(.A(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n397), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n407), .B(new_n408), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n397), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n395), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n414), .B(new_n415), .C1(new_n401), .C2(new_n402), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n418), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n406), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n313), .A2(new_n318), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n371), .B(new_n191), .C1(new_n372), .C2(new_n351), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n346), .A2(new_n353), .B1(new_n362), .B2(new_n359), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n191), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n203), .A2(G224), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  XOR2_X1   g247(.A(G116), .B(G119), .Z(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT2), .B(G113), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n357), .A3(new_n365), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT5), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n440));
  INV_X1    g254(.A(G119), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n440), .A3(new_n441), .A4(G116), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(G113), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n434), .A2(new_n435), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n399), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n433), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n437), .A2(KEYINPUT86), .A3(new_n448), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n437), .A2(new_n448), .A3(new_n433), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n451), .A2(new_n452), .B1(KEYINPUT6), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n432), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n447), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n374), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n433), .B(KEYINPUT8), .ZN(new_n464));
  INV_X1    g278(.A(new_n429), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n430), .A2(KEYINPUT7), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n429), .A2(new_n466), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n455), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n458), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G210), .B1(G237), .B2(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(KEYINPUT88), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n457), .A2(new_n458), .A3(new_n471), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n457), .A2(new_n471), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT89), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n187), .B1(new_n426), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n202), .A2(new_n203), .A3(G210), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT26), .B(G101), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n381), .A2(G134), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n209), .B1(new_n489), .B2(new_n383), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n382), .A2(new_n383), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n491), .A2(KEYINPUT67), .A3(new_n209), .A4(new_n380), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n386), .A2(new_n387), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n428), .A2(new_n390), .B1(new_n494), .B2(new_n398), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n436), .B1(new_n495), .B2(KEYINPUT30), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n428), .A2(new_n390), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n370), .A3(new_n373), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT30), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT70), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n497), .A2(new_n498), .A3(new_n501), .A4(KEYINPUT30), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n436), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n488), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(KEYINPUT28), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n497), .A2(new_n498), .A3(new_n510), .A4(new_n504), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n504), .B2(new_n495), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n507), .B(new_n508), .C1(new_n488), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n497), .A2(new_n498), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n436), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT29), .A4(new_n487), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n517), .B2(KEYINPUT75), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n514), .B(new_n518), .C1(KEYINPUT75), .C2(new_n517), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n500), .A2(new_n502), .ZN(new_n522));
  INV_X1    g336(.A(new_n496), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n505), .A2(new_n487), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT72), .B1(new_n503), .B2(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT31), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n532), .B1(new_n513), .B2(new_n488), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n521), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n519), .A2(G472), .B1(new_n534), .B2(KEYINPUT32), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n520), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT74), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n534), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n425), .A2(new_n318), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT95), .A3(new_n480), .A4(new_n313), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n270), .A2(new_n272), .A3(G119), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n269), .A2(G119), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT24), .B(G110), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT23), .B1(new_n269), .B2(G119), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n547), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT23), .A4(G119), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n198), .A2(new_n200), .A3(G146), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n222), .B1(new_n236), .B2(new_n238), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n549), .A2(new_n550), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n555), .A3(new_n552), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(new_n222), .B2(new_n212), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n201), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n201), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT22), .B(G137), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n568), .B(new_n569), .Z(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n560), .B(new_n570), .C1(new_n565), .C2(new_n566), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n294), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n572), .A2(new_n294), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n288), .B1(G234), .B2(new_n294), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n573), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n581), .A2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(KEYINPUT80), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT80), .ZN(new_n589));
  INV_X1    g403(.A(new_n581), .ZN(new_n590));
  INV_X1    g404(.A(new_n579), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n574), .B2(new_n575), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n589), .B1(new_n593), .B2(new_n586), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n482), .A2(new_n543), .A3(new_n545), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n418), .B1(new_n417), .B2(new_n294), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(KEYINPUT83), .B1(new_n423), .B2(new_n418), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n315), .B1(new_n600), .B2(new_n419), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n594), .A3(new_n588), .ZN(new_n602));
  INV_X1    g416(.A(G472), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n530), .B2(new_n533), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n537), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n598), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n536), .A2(new_n294), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n534), .B1(new_n607), .B2(G472), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n608), .A4(new_n601), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n293), .A2(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n291), .A2(new_n612), .A3(new_n292), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G478), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n299), .A2(new_n296), .ZN(new_n615));
  NAND2_X1  g429(.A1(G478), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n257), .B2(new_n312), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n451), .A2(new_n452), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n431), .B1(new_n621), .B2(new_n453), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n463), .A2(new_n464), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n465), .A2(new_n467), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n455), .A4(new_n469), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n294), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n474), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n317), .B1(new_n627), .B2(new_n478), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n306), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n610), .A2(new_n618), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n256), .A2(new_n251), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n312), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n298), .A2(new_n300), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n610), .A2(new_n629), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  OR3_X1    g454(.A1(new_n567), .A2(KEYINPUT36), .A3(new_n571), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n567), .B1(KEYINPUT36), .B2(new_n571), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n585), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n580), .B2(new_n581), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n605), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n482), .A2(new_n545), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT97), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  OAI21_X1  g464(.A(new_n628), .B1(new_n593), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n425), .A2(new_n314), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n302), .B1(new_n305), .B2(G900), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n633), .A2(new_n635), .A3(new_n312), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n543), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT98), .B(G128), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G30));
  XNOR2_X1  g472(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n480), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n257), .A2(new_n312), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n660), .A2(new_n662), .A3(new_n636), .A4(new_n317), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n582), .B1(new_n585), .B2(new_n643), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n537), .A2(KEYINPUT74), .A3(new_n539), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n541), .B1(new_n534), .B2(new_n538), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n528), .A2(new_n529), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n487), .B1(new_n516), .B2(new_n505), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n294), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n534), .A2(KEYINPUT32), .B1(new_n670), .B2(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n664), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n653), .B(KEYINPUT39), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n652), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  NAND2_X1  g495(.A1(new_n618), .A2(new_n653), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n651), .A3(new_n652), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n543), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  NAND2_X1  g499(.A1(new_n588), .A2(new_n594), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n667), .B2(new_n535), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n629), .A2(new_n618), .ZN(new_n688));
  INV_X1    g502(.A(new_n423), .ZN(new_n689));
  AND2_X1   g503(.A1(KEYINPUT101), .A2(G469), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n314), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND2_X1  g511(.A1(new_n629), .A2(new_n637), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n687), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NAND2_X1  g515(.A1(new_n664), .A2(new_n313), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n691), .A2(new_n628), .A3(new_n314), .A4(new_n692), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n543), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  AOI21_X1  g520(.A(new_n487), .B1(new_n512), .B2(new_n516), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n532), .B2(new_n531), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n530), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n520), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT102), .B(G472), .Z(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n604), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n582), .A2(new_n587), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n661), .A2(new_n306), .A3(new_n635), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n703), .A2(new_n682), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n521), .B1(new_n530), .B2(new_n708), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n607), .B2(new_n711), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n723), .B2(new_n664), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n712), .B1(new_n536), .B2(new_n294), .ZN(new_n725));
  NOR4_X1   g539(.A1(new_n725), .A2(new_n645), .A3(KEYINPUT103), .A4(new_n722), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n720), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(new_n682), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n480), .A2(new_n317), .ZN(new_n730));
  INV_X1    g544(.A(new_n424), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n408), .B(KEYINPUT104), .Z(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n417), .B2(new_n418), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n314), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n729), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n687), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n736), .A2(new_n739), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n534), .A2(KEYINPUT32), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n714), .B1(new_n535), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  INV_X1    g560(.A(new_n317), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n481), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n734), .A3(new_n654), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n687), .A2(new_n749), .A3(KEYINPUT105), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT105), .B1(new_n687), .B2(new_n749), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n276), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n418), .B1(new_n417), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n405), .A2(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n732), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT107), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n731), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n314), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n766), .A2(KEYINPUT108), .A3(new_n677), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT108), .B1(new_n766), .B2(new_n677), .ZN(new_n768));
  INV_X1    g582(.A(new_n617), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n662), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT43), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n605), .A3(new_n664), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n748), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n767), .A2(new_n768), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NAND3_X1  g591(.A1(new_n729), .A2(new_n686), .A3(new_n730), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n314), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n543), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n188), .ZN(G42));
  NAND2_X1  g597(.A1(new_n691), .A2(new_n692), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT49), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n318), .B1(new_n784), .B2(KEYINPUT49), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n714), .A4(new_n770), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n671), .B1(new_n540), .B2(new_n542), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n789), .A3(new_n660), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n543), .A2(new_n704), .B1(new_n715), .B2(new_n717), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n695), .A2(new_n700), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n695), .A2(new_n700), .A3(new_n792), .A4(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n635), .B(KEYINPUT110), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n618), .B1(new_n662), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n480), .A2(new_n306), .A3(new_n747), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n606), .A2(new_n609), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n596), .A3(new_n647), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT103), .B1(new_n713), .B2(new_n645), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n723), .A2(new_n721), .A3(new_n664), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n737), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n737), .A2(new_n807), .A3(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n752), .ZN(new_n812));
  INV_X1    g626(.A(new_n653), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n798), .A2(new_n634), .A3(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n601), .A2(new_n814), .A3(new_n664), .A4(new_n730), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n812), .A2(new_n750), .B1(new_n543), .B2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n745), .A2(new_n797), .A3(new_n811), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n661), .A2(new_n628), .A3(new_n635), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n734), .A3(new_n813), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n788), .A2(new_n645), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n727), .A2(new_n821), .A3(new_n656), .A4(new_n684), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n807), .A2(new_n720), .B1(new_n543), .B2(new_n655), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n672), .A2(new_n820), .B1(new_n543), .B2(new_n683), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n797), .A2(new_n811), .A3(new_n745), .A4(new_n816), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n818), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n823), .A2(new_n834), .A3(new_n827), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n823), .B2(new_n827), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n837), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n832), .B2(KEYINPUT113), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n791), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n748), .A2(new_n302), .A3(new_n693), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n771), .A2(new_n807), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n789), .A2(new_n842), .A3(new_n595), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n662), .A2(new_n617), .ZN(new_n845));
  INV_X1    g659(.A(new_n302), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n771), .A2(new_n846), .A3(new_n715), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n747), .B(new_n693), .C1(KEYINPUT117), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n660), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n853));
  OAI221_X1 g667(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n315), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n780), .A2(new_n781), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n847), .A2(new_n730), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n855), .B(KEYINPUT51), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n771), .A2(new_n743), .A3(new_n842), .ZN(new_n865));
  NOR2_X1   g679(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n771), .A2(new_n846), .A3(new_n715), .ZN(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n869));
  OAI221_X1 g683(.A(new_n867), .B1(new_n703), .B2(new_n868), .C1(new_n865), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n618), .ZN(new_n871));
  OAI211_X1 g685(.A(G952), .B(new_n203), .C1(new_n844), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n859), .A2(new_n862), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n855), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n864), .B(new_n873), .C1(new_n875), .C2(KEYINPUT51), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n838), .B1(new_n837), .B2(new_n829), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n811), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n878));
  INV_X1    g692(.A(new_n745), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n793), .A3(new_n838), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n482), .B(new_n545), .C1(new_n687), .C2(new_n646), .ZN(new_n882));
  INV_X1    g696(.A(new_n810), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n802), .B(new_n882), .C1(new_n883), .C2(new_n808), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n815), .A2(new_n543), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n751), .B2(new_n752), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n881), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n828), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n878), .A2(new_n880), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n877), .A2(new_n791), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n841), .A2(new_n876), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n790), .B1(new_n892), .B2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n203), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n836), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n823), .A2(new_n827), .A3(new_n834), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n817), .B2(new_n899), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n888), .A2(new_n878), .A3(new_n880), .A4(new_n887), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n294), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT56), .B1(new_n903), .B2(G210), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n454), .A2(new_n456), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n431), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n457), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n896), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n904), .B2(new_n909), .ZN(G51));
  NAND2_X1  g725(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n877), .A2(new_n913), .A3(new_n791), .A4(new_n889), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n900), .B2(new_n901), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n732), .B(KEYINPUT120), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT57), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n421), .A2(new_n422), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n902), .A2(new_n294), .A3(new_n760), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n895), .B1(new_n924), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  INV_X1    g742(.A(new_n248), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n895), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n928), .A2(new_n927), .A3(new_n929), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G60));
  AND2_X1   g748(.A1(new_n611), .A2(new_n613), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n616), .B(KEYINPUT59), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n916), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n896), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n841), .B2(new_n891), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n935), .ZN(G63));
  XNOR2_X1  g755(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n942));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n902), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n895), .B1(new_n945), .B2(new_n583), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n902), .A2(new_n944), .ZN(new_n947));
  INV_X1    g761(.A(new_n643), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n902), .A2(new_n950), .A3(new_n643), .A4(new_n944), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n946), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n946), .B(KEYINPUT61), .C1(new_n949), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n303), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n803), .B1(new_n795), .B2(new_n796), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n905), .B1(G898), .B2(new_n203), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT126), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  INV_X1    g777(.A(new_n819), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n767), .A2(new_n743), .A3(new_n768), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n824), .A2(new_n684), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n782), .A2(new_n879), .A3(new_n753), .A4(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n966), .A2(new_n968), .A3(new_n203), .A4(new_n776), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n522), .B1(KEYINPUT30), .B2(new_n495), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n217), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(G900), .B2(G953), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n799), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n687), .A2(new_n678), .A3(new_n730), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n782), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n776), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n680), .A2(new_n684), .A3(new_n824), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(new_n982), .B2(new_n203), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n974), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n974), .B2(new_n983), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G72));
  NAND4_X1  g801(.A1(new_n966), .A2(new_n968), .A3(new_n776), .A4(new_n959), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n503), .A2(new_n506), .A3(new_n487), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n978), .A2(new_n980), .A3(new_n959), .A4(new_n981), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n990), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n488), .B1(new_n524), .B2(new_n505), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(new_n997), .A3(new_n896), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n833), .A2(new_n840), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n528), .A2(new_n529), .A3(new_n507), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n990), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n999), .B2(new_n1001), .ZN(G57));
endmodule


